----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 20.04.2020 11:10:44
-- Design Name: 
-- Module Name: controlador_two_sides - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--use IEEE.STD_LOGIC_ARITH.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
library UNISIM;
use UNISIM.VComponents.all;

entity controlador_two_sides is
    Port (
		clk									: in std_logic;
        clk_100                             : in std_logic;
        dedo_ss								: out std_logic;
        dedo_mosi                           : out std_logic;
        dedo_miso                           : in std_logic;
        dedo_enable							: in std_logic;
        dedo_sclk							: out std_logic;
        frame_number					    : out std_logic_vector(7 downto 0);
        ack_ram_reading                     : out std_logic;
        interno_last_frame					: out std_logic;
        ram_reading							: in std_logic;
        DEDO_DATA_WR                        : out STD_LOGIC_VECTOR(31 downto 0);
        DEDO_ADDR_WR                        : out STD_LOGIC_VECTOR(6 downto 0);
        ROW_COLUMN                          : out STD_LOGIC_VECTOR(6 downto 0);
        START_OUT                           : out STD_LOGIC;
        enable_frame_number                 : out STD_LOGIC;
        t_ready_FIR                         : in STD_LOGIC;
        t_valid_FIR                         : out std_logic;
        r_reg_out                           : out std_logic_vector(15 downto 0)
     );
end controlador_two_sides;

architecture Behavioral of controlador_two_sides is

    -- DECLARACI�N DE SE�ALES Y TIPOS --
	type state_type is (st1_idle, st2_send_command_pause, st2_send_command, st3_send_tactel_inicial, 
								st4_send_tactel_final, st5_store_tactels, st7_interno_current_frame_update);
								
	type state_type_FIR is (st1_FIR, st2_FIR);
    
    signal state, next_state                : state_type;
    signal state_FIR, next_state_FIR        : state_type_FIR;
    signal reg_command				        : std_logic_vector(7 downto 0)  := "00000000";
	signal reg_tactel_inicial		        : std_logic_vector(7 downto 0)  := "00000000";
    signal reg_tactel_final                 : std_logic_vector(7 downto 0)  := "00000000";    
    signal byte_counter			            : std_logic_vector(2 downto 0)  := "000";
    signal contador_pausa				    : std_logic_vector(18 downto 0) := "0000000000000000000";
    signal tactel_counter		            : std_logic_vector(4 downto 0)  := "00000";
    signal row                              : std_logic_vector(2 downto 0)  := "000";
    signal column				            : std_logic_vector(3 downto 0)  := "0000";
    signal column_ret_1			            : std_logic_vector(3 downto 0)  := "0000";
    signal column_ret_2			            : std_logic_vector(3 downto 0)  := "0000";
    signal interno_current_frame		    : std_logic := '0';
    signal externo_current_frame            : std_logic := '0';
    signal pulso                            : std_logic := '0';
    signal int_dedo_addr_wr                 : std_logic_vector(7 downto 0)  := (others => '0');
    signal int_dedo_data_wr                 : std_logic_vector(31 downto 0) := (others => '0');
    signal int_frame_number    		        : std_logic_vector(7 downto 0);
    signal frame_number_stage1              : std_logic_vector(7 downto 0) := (others => '0');
    
    -- SE�AL DE START
    signal temporal_start                   : std_logic := '0';
    signal contador_start                   : integer range 0 to 4168000 := 0;
    signal duty                             : std_logic_vector(6 downto 0) := "0001010";                -- Modulaci�n de se�al para start_out
    
    -- FIR - CIRCUITO PULSO
    signal CE_DAT_REG                       : std_logic := '0';
    signal CE_RET_1                         : std_logic := '0';
    signal CE_RET_2                         : std_logic := '0';
    signal CE_PULSO_100                     : std_logic := '0';
    
    -- FIR - REGISTROS DATA Y COL-FILE
    signal data_tactel_register             : std_logic_vector(31 downto 0) := (others => '0');
    signal address_tactel_register          : std_logic_vector(6 downto 0) := (others => '0');  
    
    signal aux_addr_tactel_register         : std_logic_vector(6 downto 0) := (others => '0');
    signal aux_addr_tactel_register_slow    : std_logic_vector(6 downto 0) := (others => '0');            
          
              
    -- SPI
    signal int_dedo_ss					    : std_logic;
    signal int_dedo_mosi                    : std_logic;
    signal tactel				            : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
        
    -- ONE TACTEL
    signal contador_one_tactel              : std_logic_vector(4 downto 0) := (others => '0');
    
    -- DEPURACI�N -> BANCO DE REGISTROS
    --type t_reg_datos is array (127 downto 0) of unsigned(31 downto 0);
--    type t_reg_datos is array (0 to 1023) of natural;
--    type t_reg_datos is array (0 to 1023) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (98, 1328, 3672, 6741, 10032, 13017, 15245, 16421, 16461, 15501, 13873, 12037, 10492, 9678, 9893, 11232, 13568, 16569, 19764, 22625, 24666, 25533, 25070, 23345, 20643, 17409, 14169, 11431, 9592, 8866, 9251, 10524, 12295, 14075, 15378, 15812, 15153, 13397, 10757, 7628, 4516, 1943, 352, 25, 1028, 3201, 6188, 9499, 12605, 15031, 16445, 16719, 15944, 14418, 12582, 10935, 9936, 9918, 11019, 13156, 16036, 19210, 22154, 24366, 25460, 25237, 23722, 21159, 17967, 14665, 11771, 9712, 8746, 8911, 10029, 11737, 13559, 15001, 15644, 15226, 13697, 11228, 8182, 5048, 2355, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590, 15430, 15250, 13955, 11671, 8727, 5593, 2798, 566, 0, 770, 2758, 5643, 8954, 12162, 14773, 16421, 16932, 16356, 14951, 13136, 11406, 10236, 9991, 10851, 12779, 15520, 18652, 21659, 24026, 25340, 25358, 24062, 21654, 18525, 15180, 12148, 9880, 8673, 8611, 9558, 11183, 13027, 14590);
    
--    type t_reg_datos is array (0 to 2047) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (20281, 19442, 16957, 15142, 15412, 15158, 15446, 15015, 15796, 13576, 13213, 14746, 14148, 13681, 14541, 16329, 16067, 17112, 17673, 17879, 17338, 16618, 17513, 17677, 18974, 19412, 19299, 20713, 20716, 21630, 19675, 17264, 17171, 15561, 14850, 14784, 14268, 13055, 12547, 12652, 15122, 16961, 15195, 15539, 15896, 16354, 18070, 17031, 15867, 16308, 15920, 16433, 15532, 18360, 21149, 20358, 20118, 20773, 18637, 15919, 16950, 15582, 14798, 14490, 13714, 12949, 12545, 12596, 14971, 15943, 14995, 15356, 15244, 15672, 15149, 16057, 12456, 12160, 14705, 14746, 17536, 19683, 20632, 19339, 18951, 18961, 18166, 16160, 14775, 13998, 13819, 14098, 13968, 14087, 13927, 14190, 13695, 15172, 15826, 15349, 15793, 15411, 15282, 15425, 13628, 10017, 13746, 17765, 18410, 19097, 18160, 18291, 18266, 18194, 16299, 14385, 14564, 14430, 14794, 15266, 14333, 13756, 13479, 13309, 14106, 14906, 15300, 15144, 15461, 16010, 15456, 16309, 13637, 10992, 11725, 11282, 11449, 11483, 11226, 11807, 10600, 14305, 16406, 15236, 13275, 13058, 15040, 13489, 14385, 13898, 13520, 14624, 14786, 15443, 16125, 15897, 16159, 16090, 16773, 16294, 17475, 13735, 13670, 18340, 18214, 19152, 18688, 18990, 19240, 18986, 18450, 16352, 15067, 14897, 14771, 13998, 13388, 13457, 13339, 13298, 13285, 13327, 13245, 13388, 13092, 14315, 16772, 14728, 11917, 10636, 15085, 21140, 22611, 22406, 19945, 18489, 18989, 17788, 16992, 14503, 12555, 13098, 12361, 12425, 12993, 13356, 13007, 12966, 16652, 20103, 14402, 12960, 15909, 16334, 17999, 14797, 12790, 12737, 15005, 21705, 24848, 24482, 20347, 18059, 18770, 18263, 18819, 18002, 19501, 14603, 9666, 13565, 13866, 12085, 13051, 17623, 19252, 14209, 14067, 15731, 15216, 18963, 15817, 11225, 14981, 17980, 20281, 24541, 22807, 20467, 19093, 17833, 17734, 17626, 14109, 11981, 12690, 12902, 14158, 12030, 12482, 11230, 12450, 15248, 18058, 13732, 10762, 13912, 12626, 13377, 12833, 13384, 12527, 15303, 19022, 17438, 14309, 12046, 12024, 11579, 10825, 10179, 9118, 8125, 2635, 0, 255, 65, 1114, 3226, 7181, 4937, 4904, 5229, 2274, 2739, 3468, 3943, 3801, 7301, 6678, 7174, 10900, 8869, 8498, 8904, 9335, 9643, 7035, 3477, 966, 593, 639, 616, 637, 614, 646, 432, 0, 920, 1607, 2215, 1551, 3975, 8143, 8214, 10267, 9741, 7938, 10131, 10187, 7457, 5714, 6561, 8137, 8270, 7601, 2265, 0, 225, 0, 67, 0, 14, 0, 26, 0, 137, 0, 490, 0, 3741, 7569, 6772, 8447, 7694, 8055, 7896, 7942, 7960, 7852, 8708, 10921, 4059, 0, 455, 0, 149, 0, 108, 0, 273, 0, 1795, 1923, 0, 581, 0, 2464, 5584, 6427, 7625, 6219, 6980, 7178, 7515, 9055, 9759, 8363, 8337, 3322, 0, 396, 0, 113, 0, 22, 0, 0, 5, 0, 25, 0, 85, 0, 1129, 5119, 7333, 7720, 7425, 6328, 7226, 7642, 8519, 10360, 9287, 10455, 4203, 0, 502, 0, 146, 0, 29, 0, 0, 0, 0, 22, 0, 107, 0, 365, 0, 3117, 7916, 6425, 6725, 6224, 6632, 7095, 7462, 9068, 9327, 9414, 9186, 9628, 8807, 10461, 4833, 0, 1652, 748, 0, 56, 0, 0, 79, 0, 1299, 5605, 7450, 7420, 8089, 7137, 7347, 7928, 7175, 8053, 8066, 7902, 6757, 1869, 0, 216, 0, 165, 0, 1621, 6307, 2332, 684, 2183, 0, 958, 48, 3849, 7098, 6110, 6637, 6305, 6562, 6266, 7096, 8173, 7923, 8830, 8909, 8653, 7891, 6772, 2250, 0, 0, 1635, 7379, 8126, 8533, 10605, 7486, 1583, 3259, 5942, 7265, 9388, 10075, 10243, 10946, 13124, 15126, 11046, 7483, 9598, 10056, 10725, 9051, 7840, 7345, 7244, 6372, 3654, 2900, 3028, 2991, 2975, 3060, 2833, 3762, 6458, 10692, 11310, 10331, 10642, 12155, 15508, 15761, 16054, 13437, 11339, 14072, 13996, 13475, 12873, 11615, 12032, 12772, 10522, 7813, 8735, 8864, 8034, 11356, 15652, 11520, 7766, 9196, 10968, 13339, 11543, 9800, 11402, 15953, 17335, 17562, 17249, 15480, 16118, 15775, 15985, 15834, 16004, 15238, 12837, 13847, 12237, 10779, 9816, 11283, 14596, 15024, 13224, 8358, 11357, 13157, 13102, 14028, 11838, 15129, 18273, 18704, 20247, 19379, 17872, 16548, 16950, 16816, 14881, 15317, 15546, 15735, 14612, 14881, 14038, 11290, 11287, 13466, 14409, 16901, 14288, 10132, 11380, 10918, 10863, 11461, 9962, 15185, 20963, 20440, 20258, 19894, 19252, 16721, 17812, 14863, 14061, 16449, 16516, 15066, 13806, 13506, 10511, 11441, 14931, 16351, 18347, 16891, 14023, 17214, 17828, 17517, 14797, 11401, 17224, 20947, 20630, 21565, 21323, 20805, 20329, 19229, 16600, 14057, 14093, 14225, 14196, 14227, 14176, 14268, 14082, 14738, 16248, 17976, 16379, 13947, 16160, 16820, 17745, 15421, 9689, 14072, 19190, 19611, 20900, 20795, 20884, 20767, 19269, 18155, 15030, 13536, 14480, 14349, 14608, 14567, 15113, 14789, 13605, 15000, 18023, 18708, 18917, 16311, 16784, 19585, 18798, 20182, 16139, 12803, 13937, 13105, 14026, 12562, 17046, 21469, 18214, 15494, 14608, 14335, 15595, 15708, 14321, 15321, 15338, 14314, 14613, 17024, 18941, 18795, 16204, 16422, 19190, 18850, 20022, 15168, 11334, 17152, 19513, 19939, 21029, 20792, 20773, 20717, 17569, 16641, 16440, 16247, 16519, 16473, 15031, 14039, 14823, 14592, 14811, 14553, 14947, 14206, 16551, 18821, 19041, 18723, 14112, 11088, 15502, 19163, 18715, 19994, 20587, 20987, 19883, 17590, 16950, 15847, 14356, 15459, 16560, 15901, 15070, 13276, 11730, 13861, 15860, 17149, 18856, 18175, 17988, 18517, 18748, 19746, 14428, 10815, 16516, 19356, 19377, 19850, 19812, 19905, 19801, 19949, 19712, 20165, 18572, 16401, 17048, 14936, 15206, 15173, 14653, 16057, 17998, 18218, 15804, 16545, 18333, 18704, 19847, 15051, 9722, 16100, 19637, 19678, 20378, 19918, 20081, 19661, 18705, 16859, 15487, 14896, 14466, 14827, 15808, 15330, 17227, 14345, 13736, 17507, 17594, 18899, 18851, 18930, 18910, 18884, 18956, 18811, 19247, 19599, 20003, 20339, 20718, 20920, 20182, 19225, 17674, 17306, 17460, 17100, 16879, 16271, 16435, 16475, 16062, 16113, 17085, 18384, 20138, 21258, 20815, 20745, 19765, 21504, 18647, 15977, 18963, 20229, 21507, 22091, 22165, 21312, 20594, 20249, 20086, 18347, 17225, 17521, 17407, 17412, 17514, 17241, 18278, 19862, 20198, 21729, 23169, 23408, 22883, 21507, 22092, 22299, 21487, 20842, 20550, 21584, 21844, 21899, 21064, 20738, 20364, 18778, 17499, 17717, 17025, 16836, 16756, 16831, 17719, 16325, 15754, 16647, 16994, 18597, 19550, 18348, 18831, 18222, 20358, 15940, 11093, 12523, 11935, 12015, 12410, 11312, 15033, 17790, 16113, 16788, 13767, 13143, 15471, 15399, 15222, 14088, 12380, 10638, 13166, 15917, 16319, 17270, 16409, 16357, 15903, 18089, 13695, 11388, 11669, 13521, 17531, 18329, 17603, 16121, 17036, 15898, 16002, 13961, 12099, 13014, 14431, 14699, 15430, 13642, 11681, 12209, 12095, 11880, 12510, 11113, 15743, 20361, 20093, 19120, 17094, 20220, 20611, 19873, 20153, 20818, 20987, 20723, 20660, 18043, 16835, 16638, 17312, 18536, 18256, 18722, 18593, 18417, 18077, 19014, 20006, 20503, 21940, 21918, 21666, 21331, 21651, 21623, 20151, 20580, 20505, 19919, 19328, 19539, 20230, 19988, 20130, 20013, 20156, 19934, 20203, 17684, 16194, 16945, 17566, 16462, 16662, 18657, 19169, 20838, 20501, 20893, 20445, 20656, 20855, 19221, 19501, 19071, 18286, 17645, 18226, 19728, 19857, 20516, 19829, 17174, 15080, 15992, 16471, 15062, 14414, 13557, 13869, 14218, 15119, 17115, 18691, 18914, 18580, 18709, 18616, 18724, 18551, 18863, 18133, 18364, 15830, 13589, 15120, 14713, 15246, 16053, 15521, 15152, 15590, 15633, 15438, 15363, 14548, 13330, 13065, 14661, 15036, 17719, 18408, 18015, 20394, 20470, 21159, 20305, 19571, 19192, 19492, 19246, 16803, 17856, 18577, 18772, 18754, 18662, 19031, 18623, 19072, 18914, 18941, 19025, 18804, 19273, 17786, 16972, 18806, 19569, 20623, 20650, 19968, 19779, 18803, 18441, 17596, 18267, 19323, 17268, 17503, 18558, 18968, 20062, 19570, 19947, 19936, 20530, 20483, 18232, 17304, 16281, 16731, 17839, 19169, 17754, 18701, 19890, 21362, 20445, 19595, 20930, 19705, 20613, 20545, 20641, 20571, 20645, 20532, 20743, 20109, 20049, 21585, 21041, 21547, 20597, 19792, 19844, 18925, 18633, 19976, 20369, 18756, 19835, 20773, 22396, 21882, 21399, 22636, 21728, 21979, 22119, 21897, 22238, 21543, 20891, 20668, 20976, 21683, 21640, 21151, 22192, 21458, 19742, 20137, 19120, 18131, 18930, 19300, 19174, 19329, 19066, 19537, 18628, 21372, 22940, 22010, 23210, 22055, 23772, 24015, 22753, 22965, 22504, 22424, 22446, 22208, 22751, 22751, 22768, 21805, 21795, 21022, 19172, 20004, 20124, 21045, 22316, 21595, 20749, 20764, 22691, 23159, 21718, 21988, 23110, 22205, 23220, 24502, 23425, 24121, 23879, 23631, 23717, 23640, 23736, 23589, 23865, 22931, 21683, 21929, 22501, 21997, 21229, 22531, 23140, 22670, 22846, 22199, 22367, 21840, 21632, 22843, 23079, 22151, 22119, 23459, 23930, 24182, 22964, 22752, 22965, 22415, 23357, 23692, 22440, 22035, 21641, 21550, 22266, 22083, 22797, 23654, 23153, 22047, 22150, 22662, 22496, 22577, 22540, 22546, 22567, 22583, 23494, 24453, 24971, 23851, 23081, 23220, 22914, 22993, 22507, 22303, 22661, 22018, 21586, 22611, 21584, 23130, 24542, 22856, 22155, 22283, 22374, 23379, 22852, 22123, 23380, 22802, 23146, 23936, 24669, 25235, 24608, 24078, 23536, 22986, 22137, 21445, 22548, 23201, 23025, 23122, 23049, 23124, 23024, 23173, 22101, 20162, 20176, 21106, 21454, 21176, 21326, 21634, 21672, 22184, 22296, 23203, 23916, 23891, 22567, 21314, 20336, 20060, 20993, 21167, 21249, 21164, 21288, 20632, 20546, 20042, 21467, 23147, 21406, 19880, 19827, 20252, 21058, 20462, 19998, 21131, 20520, 19988, 20137, 20057, 20108, 20072, 20112, 19919, 19052, 18484, 18284, 18523, 18777, 17661, 17295, 16575, 17365, 18433, 20520, 20103, 17864, 18706, 19168, 20000, 20184, 19944, 19534, 18360, 19710, 21108, 21214, 22027, 21600, 21043, 19431, 18358, 17862, 17880, 17746, 17216, 17310, 16892, 16206, 16297, 16576, 16563, 16549, 16614, 16468, 16755, 16172, 17987, 19090, 18354, 18165, 19711, 19827, 18805, 20217, 19896, 18950, 18080, 17749, 17409, 17081, 16151, 15824, 14641, 14602, 15526, 15361, 14517, 15111, 14635, 16489, 17884, 16678, 17309, 17983, 19085, 18465, 18285, 17317, 18171, 18945, 18097, 19197, 19909, 19158, 18823, 18776, 19008, 18520, 19528, 16160, 12615, 13650, 13447, 14573, 14711, 14870, 16331, 16913, 16365, 16170, 17020, 18034, 17324, 16363, 15948, 17105, 18052, 18041, 18207, 18521, 17600, 16925, 16203, 15367, 15007, 14359, 14672, 14163, 13598, 13649, 13702, 14018, 14805, 14622, 14979, 15816, 15701, 16476, 17066, 16907, 16963, 16981, 16876, 17154, 17083, 18845, 19087, 17665, 18386, 16635, 15991, 14861, 14353, 15129, 14246, 14322, 13996, 14161, 14402, 14842, 14656, 14770, 15819, 15910, 16360, 15903, 16336, 15398, 11657, 14541, 18052, 17135, 17478, 17790, 18248, 17843, 17523, 16147, 15325, 13228, 11507, 13367, 13622, 13703, 13553, 13815, 13306, 14774, 14717, 12966, 13157, 14140, 15909, 16019, 16663, 13971, 15076, 18813, 18232, 19076, 18629, 17955, 17800, 17424, 17025, 15942, 15830, 15862, 15995, 15034, 14499, 14539, 14189, 14973, 15755, 14871, 12697, 12235, 12300, 13476, 15618, 15720, 16529, 14521, 15926, 18815, 17862, 18357, 18067, 18263, 18083, 18275, 17001, 15817, 14654, 13660, 14348, 13337, 14686, 12378, 12461, 15777, 15419, 13850, 13204, 14400, 14703, 16901, 17308, 14988, 12878, 16271, 18966, 18395, 19010, 18285, 17857, 17803, 17834, 18601, 17024, 15687, 16041, 16588, 16871, 15002, 14425, 14693, 15134, 15743, 15512, 15672, 15517, 15720, 15354, 16740, 18778, 15919, 16679, 19339, 18116, 17912, 18139, 17935, 17791, 17812, 18008, 16714, 15010, 16251, 16784, 16585, 15701, 15116, 14448, 15071, 16740, 17171, 17107, 16663, 17124, 17614, 18261, 18404, 18764, 18443, 18376, 19021, 17875, 17218, 17698, 17424, 17199, 17121, 17164, 17100, 17214, 17007, 17419, 16079, 14938, 16210, 16952, 17556, 16829, 15975, 16347, 17029, 17410, 17629, 18323, 18434, 18004, 18807, 18448, 17900, 18317, 18301, 18236, 17581, 18060, 17616, 16960, 17066, 17034, 16113, 15246, 15743, 16570, 15383, 15784, 17132, 16029, 16049, 16903, 17405, 17475, 17765, 17661, 17717, 17680, 17716, 17660, 17860, 18320, 18572, 18097, 18032, 17589, 15921, 14980, 15054, 15033, 15140, 16526, 13353, 10618, 15439, 16819, 16681, 16398, 15656, 16736, 16983, 17792, 19086, 17095, 16842, 18838, 17748, 17796, 17886, 18139, 18496, 18178, 18269, 17407, 16940, 17342, 17239, 15912, 14954, 15222, 15109, 15136, 15184, 15029, 15598, 16415, 17089, 17636, 18048, 18791, 17820, 17721, 18177, 17058, 16788, 17769, 18406, 18055, 17898, 16939, 16416, 15497, 13603, 14502, 14278, 15185, 14619, 13733, 15205, 15537, 16479, 15931, 15313, 16704, 17438, 17835, 17097, 15877, 14594, 16431, 18264, 17037, 17322, 17181, 17167, 17351, 16930, 17808, 15045, 12894, 12793, 13546, 14110, 12176, 10790, 13836, 17425, 15847, 15136, 13414, 13862, 14867, 15067, 16260, 16048, 14548, 16361, 18112, 17303, 17213, 17507, 17628, 17411, 17414, 16276, 16212, 15062, 13954, 12458, 12290, 12812, 10822, 13126, 16335, 17302, 15525, 14296, 14607, 14526, 14441, 14723, 14086, 16224, 18269, 17334, 17375, 17076, 17724, 17604, 17275, 17266, 17348, 15843, 13985, 15081, 14478, 14844, 13655, 13911, 16738, 16893, 17977, 16885, 15335, 16273, 16740, 17285, 18492, 18491, 18002, 18105, 18475, 18117, 17811, 17633, 17935, 17581, 17696, 16669, 16406, 17296, 16970, 17139, 17051, 17086, 17081, 17209, 18090, 16558, 14379, 13579, 15512, 17210, 17202, 14957, 15364, 18369, 18080, 18562, 18350, 18228, 18611, 18019, 17835, 17374, 16867, 16650, 15941, 16107, 16678, 16272, 16083, 15410, 16690, 17332, 16519, 15884, 15363, 15054, 16548, 17279, 16660, 15713, 16437, 18564, 17841, 18216, 17994, 18153, 17990, 18223, 17192, 16175, 16085, 16095, 16032, 16423, 16627, 16036, 15876, 16265, 16877, 16682, 16139, 16147, 16167, 17701, 18223, 17249, 18594, 19373, 19811, 19952, 19605, 19665, 18873, 18260, 17844, 18564, 17596, 16249, 16597, 16242, 16554, 16483, 15998, 15924, 15965, 15802, 15844, 15857, 15783, 15947, 15608, 16681, 17591, 17964, 19396, 19880, 19763, 19132, 19458, 19256, 17883, 17782, 18291, 17106, 15893, 17079, 17446, 17765, 17078, 16026, 15909, 16355, 17300, 17428, 16956, 17340, 18382, 18010, 18212, 18405, 18846, 19310, 19805, 19449, 19257, 18809, 18539, 18562, 17917, 17967, 17933, 17914, 17995, 17824, 18173, 17054, 15949, 15693, 15648, 16941, 17157, 16957, 17892, 18463, 18091, 18349, 18712, 18970, 18792, 18313, 18964, 19168);

--    type t_reg_datos is array (0 to 16383) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (20281, 19442, 16957, 15142, 15412, 15158, 15446, 15015, 15796, 13576, 13213, 14746, 14148, 13681, 14541, 16329, 16067, 17112, 17673, 17879, 17338, 16618, 17513, 17677, 18974, 19412, 19299, 20713, 20716, 21630, 19675, 17264, 17171, 15561, 14850, 14784, 14268, 13055, 12547, 12652, 15122, 16961, 15195, 15539, 15896, 16354, 18070, 17031, 15867, 16308, 15920, 16433, 15532, 18360, 21149, 20358, 20118, 20773, 18637, 15919, 16950, 15582, 14798, 14490, 13714, 12949, 12545, 12596, 14971, 15943, 14995, 15356, 15244, 15672, 15149, 16057, 12456, 12160, 14705, 14746, 17536, 19683, 20632, 19339, 18951, 18961, 18166, 16160, 14775, 13998, 13819, 14098, 13968, 14087, 13927, 14190, 13695, 15172, 15826, 15349, 15793, 15411, 15282, 15425, 13628, 10017, 13746, 17765, 18410, 19097, 18160, 18291, 18266, 18194, 16299, 14385, 14564, 14430, 14794, 15266, 14333, 13756, 13479, 13309, 14106, 14906, 15300, 15144, 15461, 16010, 15456, 16309, 13637, 10992, 11725, 11282, 11449, 11483, 11226, 11807, 10600, 14305, 16406, 15236, 13275, 13058, 15040, 13489, 14385, 13898, 13520, 14624, 14786, 15443, 16125, 15897, 16159, 16090, 16773, 16294, 17475, 13735, 13670, 18340, 18214, 19152, 18688, 18990, 19240, 18986, 18450, 16352, 15067, 14897, 14771, 13998, 13388, 13457, 13339, 13298, 13285, 13327, 13245, 13388, 13092, 14315, 16772, 14728, 11917, 10636, 15085, 21140, 22611, 22406, 19945, 18489, 18989, 17788, 16992, 14503, 12555, 13098, 12361, 12425, 12993, 13356, 13007, 12966, 16652, 20103, 14402, 12960, 15909, 16334, 17999, 14797, 12790, 12737, 15005, 21705, 24848, 24482, 20347, 18059, 18770, 18263, 18819, 18002, 19501, 14603, 9666, 13565, 13866, 12085, 13051, 17623, 19252, 14209, 14067, 15731, 15216, 18963, 15817, 11225, 14981, 17980, 20281, 24541, 22807, 20467, 19093, 17833, 17734, 17626, 14109, 11981, 12690, 12902, 14158, 12030, 12482, 11230, 12450, 15248, 18058, 13732, 10762, 13912, 12626, 13377, 12833, 13384, 12527, 15303, 19022, 17438, 14309, 12046, 12024, 11579, 10825, 10179, 9118, 8125, 2635, 0, 255, 65, 1114, 3226, 7181, 4937, 4904, 5229, 2274, 2739, 3468, 3943, 3801, 7301, 6678, 7174, 10900, 8869, 8498, 8904, 9335, 9643, 7035, 3477, 966, 593, 639, 616, 637, 614, 646, 432, 0, 920, 1607, 2215, 1551, 3975, 8143, 8214, 10267, 9741, 7938, 10131, 10187, 7457, 5714, 6561, 8137, 8270, 7601, 2265, 0, 225, 0, 67, 0, 14, 0, 26, 0, 137, 0, 490, 0, 3741, 7569, 6772, 8447, 7694, 8055, 7896, 7942, 7960, 7852, 8708, 10921, 4059, 0, 455, 0, 149, 0, 108, 0, 273, 0, 1795, 1923, 0, 581, 0, 2464, 5584, 6427, 7625, 6219, 6980, 7178, 7515, 9055, 9759, 8363, 8337, 3322, 0, 396, 0, 113, 0, 22, 0, 0, 5, 0, 25, 0, 85, 0, 1129, 5119, 7333, 7720, 7425, 6328, 7226, 7642, 8519, 10360, 9287, 10455, 4203, 0, 502, 0, 146, 0, 29, 0, 0, 0, 0, 22, 0, 107, 0, 365, 0, 3117, 7916, 6425, 6725, 6224, 6632, 7095, 7462, 9068, 9327, 9414, 9186, 9628, 8807, 10461, 4833, 0, 1652, 748, 0, 56, 0, 0, 79, 0, 1299, 5605, 7450, 7420, 8089, 7137, 7347, 7928, 7175, 8053, 8066, 7902, 6757, 1869, 0, 216, 0, 165, 0, 1621, 6307, 2332, 684, 2183, 0, 958, 48, 3849, 7098, 6110, 6637, 6305, 6562, 6266, 7096, 8173, 7923, 8830, 8909, 8653, 7891, 6772, 2250, 0, 0, 1635, 7379, 8126, 8533, 10605, 7486, 1583, 3259, 5942, 7265, 9388, 10075, 10243, 10946, 13124, 15126, 11046, 7483, 9598, 10056, 10725, 9051, 7840, 7345, 7244, 6372, 3654, 2900, 3028, 2991, 2975, 3060, 2833, 3762, 6458, 10692, 11310, 10331, 10642, 12155, 15508, 15761, 16054, 13437, 11339, 14072, 13996, 13475, 12873, 11615, 12032, 12772, 10522, 7813, 8735, 8864, 8034, 11356, 15652, 11520, 7766, 9196, 10968, 13339, 11543, 9800, 11402, 15953, 17335, 17562, 17249, 15480, 16118, 15775, 15985, 15834, 16004, 15238, 12837, 13847, 12237, 10779, 9816, 11283, 14596, 15024, 13224, 8358, 11357, 13157, 13102, 14028, 11838, 15129, 18273, 18704, 20247, 19379, 17872, 16548, 16950, 16816, 14881, 15317, 15546, 15735, 14612, 14881, 14038, 11290, 11287, 13466, 14409, 16901, 14288, 10132, 11380, 10918, 10863, 11461, 9962, 15185, 20963, 20440, 20258, 19894, 19252, 16721, 17812, 14863, 14061, 16449, 16516, 15066, 13806, 13506, 10511, 11441, 14931, 16351, 18347, 16891, 14023, 17214, 17828, 17517, 14797, 11401, 17224, 20947, 20630, 21565, 21323, 20805, 20329, 19229, 16600, 14057, 14093, 14225, 14196, 14227, 14176, 14268, 14082, 14738, 16248, 17976, 16379, 13947, 16160, 16820, 17745, 15421, 9689, 14072, 19190, 19611, 20900, 20795, 20884, 20767, 19269, 18155, 15030, 13536, 14480, 14349, 14608, 14567, 15113, 14789, 13605, 15000, 18023, 18708, 18917, 16311, 16784, 19585, 18798, 20182, 16139, 12803, 13937, 13105, 14026, 12562, 17046, 21469, 18214, 15494, 14608, 14335, 15595, 15708, 14321, 15321, 15338, 14314, 14613, 17024, 18941, 18795, 16204, 16422, 19190, 18850, 20022, 15168, 11334, 17152, 19513, 19939, 21029, 20792, 20773, 20717, 17569, 16641, 16440, 16247, 16519, 16473, 15031, 14039, 14823, 14592, 14811, 14553, 14947, 14206, 16551, 18821, 19041, 18723, 14112, 11088, 15502, 19163, 18715, 19994, 20587, 20987, 19883, 17590, 16950, 15847, 14356, 15459, 16560, 15901, 15070, 13276, 11730, 13861, 15860, 17149, 18856, 18175, 17988, 18517, 18748, 19746, 14428, 10815, 16516, 19356, 19377, 19850, 19812, 19905, 19801, 19949, 19712, 20165, 18572, 16401, 17048, 14936, 15206, 15173, 14653, 16057, 17998, 18218, 15804, 16545, 18333, 18704, 19847, 15051, 9722, 16100, 19637, 19678, 20378, 19918, 20081, 19661, 18705, 16859, 15487, 14896, 14466, 14827, 15808, 15330, 17227, 14345, 13736, 17507, 17594, 18899, 18851, 18930, 18910, 18884, 18956, 18811, 19247, 19599, 20003, 20339, 20718, 20920, 20182, 19225, 17674, 17306, 17460, 17100, 16879, 16271, 16435, 16475, 16062, 16113, 17085, 18384, 20138, 21258, 20815, 20745, 19765, 21504, 18647, 15977, 18963, 20229, 21507, 22091, 22165, 21312, 20594, 20249, 20086, 18347, 17225, 17521, 17407, 17412, 17514, 17241, 18278, 19862, 20198, 21729, 23169, 23408, 22883, 21507, 22092, 22299, 21487, 20842, 20550, 21584, 21844, 21899, 21064, 20738, 20364, 18778, 17499, 17717, 17025, 16836, 16756, 16831, 17719, 16325, 15754, 16647, 16994, 18597, 19550, 18348, 18831, 18222, 20358, 15940, 11093, 12523, 11935, 12015, 12410, 11312, 15033, 17790, 16113, 16788, 13767, 13143, 15471, 15399, 15222, 14088, 12380, 10638, 13166, 15917, 16319, 17270, 16409, 16357, 15903, 18089, 13695, 11388, 11669, 13521, 17531, 18329, 17603, 16121, 17036, 15898, 16002, 13961, 12099, 13014, 14431, 14699, 15430, 13642, 11681, 12209, 12095, 11880, 12510, 11113, 15743, 20361, 20093, 19120, 17094, 20220, 20611, 19873, 20153, 20818, 20987, 20723, 20660, 18043, 16835, 16638, 17312, 18536, 18256, 18722, 18593, 18417, 18077, 19014, 20006, 20503, 21940, 21918, 21666, 21331, 21651, 21623, 20151, 20580, 20505, 19919, 19328, 19539, 20230, 19988, 20130, 20013, 20156, 19934, 20203, 17684, 16194, 16945, 17566, 16462, 16662, 18657, 19169, 20838, 20501, 20893, 20445, 20656, 20855, 19221, 19501, 19071, 18286, 17645, 18226, 19728, 19857, 20516, 19829, 17174, 15080, 15992, 16471, 15062, 14414, 13557, 13869, 14218, 15119, 17115, 18691, 18914, 18580, 18709, 18616, 18724, 18551, 18863, 18133, 18364, 15830, 13589, 15120, 14713, 15246, 16053, 15521, 15152, 15590, 15633, 15438, 15363, 14548, 13330, 13065, 14661, 15036, 17719, 18408, 18015, 20394, 20470, 21159, 20305, 19571, 19192, 19492, 19246, 16803, 17856, 18577, 18772, 18754, 18662, 19031, 18623, 19072, 18914, 18941, 19025, 18804, 19273, 17786, 16972, 18806, 19569, 20623, 20650, 19968, 19779, 18803, 18441, 17596, 18267, 19323, 17268, 17503, 18558, 18968, 20062, 19570, 19947, 19936, 20530, 20483, 18232, 17304, 16281, 16731, 17839, 19169, 17754, 18701, 19890, 21362, 20445, 19595, 20930, 19705, 20613, 20545, 20641, 20571, 20645, 20532, 20743, 20109, 20049, 21585, 21041, 21547, 20597, 19792, 19844, 18925, 18633, 19976, 20369, 18756, 19835, 20773, 22396, 21882, 21399, 22636, 21728, 21979, 22119, 21897, 22238, 21543, 20891, 20668, 20976, 21683, 21640, 21151, 22192, 21458, 19742, 20137, 19120, 18131, 18930, 19300, 19174, 19329, 19066, 19537, 18628, 21372, 22940, 22010, 23210, 22055, 23772, 24015, 22753, 22965, 22504, 22424, 22446, 22208, 22751, 22751, 22768, 21805, 21795, 21022, 19172, 20004, 20124, 21045, 22316, 21595, 20749, 20764, 22691, 23159, 21718, 21988, 23110, 22205, 23220, 24502, 23425, 24121, 23879, 23631, 23717, 23640, 23736, 23589, 23865, 22931, 21683, 21929, 22501, 21997, 21229, 22531, 23140, 22670, 22846, 22199, 22367, 21840, 21632, 22843, 23079, 22151, 22119, 23459, 23930, 24182, 22964, 22752, 22965, 22415, 23357, 23692, 22440, 22035, 21641, 21550, 22266, 22083, 22797, 23654, 23153, 22047, 22150, 22662, 22496, 22577, 22540, 22546, 22567, 22583, 23494, 24453, 24971, 23851, 23081, 23220, 22914, 22993, 22507, 22303, 22661, 22018, 21586, 22611, 21584, 23130, 24542, 22856, 22155, 22283, 22374, 23379, 22852, 22123, 23380, 22802, 23146, 23936, 24669, 25235, 24608, 24078, 23536, 22986, 22137, 21445, 22548, 23201, 23025, 23122, 23049, 23124, 23024, 23173, 22101, 20162, 20176, 21106, 21454, 21176, 21326, 21634, 21672, 22184, 22296, 23203, 23916, 23891, 22567, 21314, 20336, 20060, 20993, 21167, 21249, 21164, 21288, 20632, 20546, 20042, 21467, 23147, 21406, 19880, 19827, 20252, 21058, 20462, 19998, 21131, 20520, 19988, 20137, 20057, 20108, 20072, 20112, 19919, 19052, 18484, 18284, 18523, 18777, 17661, 17295, 16575, 17365, 18433, 20520, 20103, 17864, 18706, 19168, 20000, 20184, 19944, 19534, 18360, 19710, 21108, 21214, 22027, 21600, 21043, 19431, 18358, 17862, 17880, 17746, 17216, 17310, 16892, 16206, 16297, 16576, 16563, 16549, 16614, 16468, 16755, 16172, 17987, 19090, 18354, 18165, 19711, 19827, 18805, 20217, 19896, 18950, 18080, 17749, 17409, 17081, 16151, 15824, 14641, 14602, 15526, 15361, 14517, 15111, 14635, 16489, 17884, 16678, 17309, 17983, 19085, 18465, 18285, 17317, 18171, 18945, 18097, 19197, 19909, 19158, 18823, 18776, 19008, 18520, 19528, 16160, 12615, 13650, 13447, 14573, 14711, 14870, 16331, 16913, 16365, 16170, 17020, 18034, 17324, 16363, 15948, 17105, 18052, 18041, 18207, 18521, 17600, 16925, 16203, 15367, 15007, 14359, 14672, 14163, 13598, 13649, 13702, 14018, 14805, 14622, 14979, 15816, 15701, 16476, 17066, 16907, 16963, 16981, 16876, 17154, 17083, 18845, 19087, 17665, 18386, 16635, 15991, 14861, 14353, 15129, 14246, 14322, 13996, 14161, 14402, 14842, 14656, 14770, 15819, 15910, 16360, 15903, 16336, 15398, 11657, 14541, 18052, 17135, 17478, 17790, 18248, 17843, 17523, 16147, 15325, 13228, 11507, 13367, 13622, 13703, 13553, 13815, 13306, 14774, 14717, 12966, 13157, 14140, 15909, 16019, 16663, 13971, 15076, 18813, 18232, 19076, 18629, 17955, 17800, 17424, 17025, 15942, 15830, 15862, 15995, 15034, 14499, 14539, 14189, 14973, 15755, 14871, 12697, 12235, 12300, 13476, 15618, 15720, 16529, 14521, 15926, 18815, 17862, 18357, 18067, 18263, 18083, 18275, 17001, 15817, 14654, 13660, 14348, 13337, 14686, 12378, 12461, 15777, 15419, 13850, 13204, 14400, 14703, 16901, 17308, 14988, 12878, 16271, 18966, 18395, 19010, 18285, 17857, 17803, 17834, 18601, 17024, 15687, 16041, 16588, 16871, 15002, 14425, 14693, 15134, 15743, 15512, 15672, 15517, 15720, 15354, 16740, 18778, 15919, 16679, 19339, 18116, 17912, 18139, 17935, 17791, 17812, 18008, 16714, 15010, 16251, 16784, 16585, 15701, 15116, 14448, 15071, 16740, 17171, 17107, 16663, 17124, 17614, 18261, 18404, 18764, 18443, 18376, 19021, 17875, 17218, 17698, 17424, 17199, 17121, 17164, 17100, 17214, 17007, 17419, 16079, 14938, 16210, 16952, 17556, 16829, 15975, 16347, 17029, 17410, 17629, 18323, 18434, 18004, 18807, 18448, 17900, 18317, 18301, 18236, 17581, 18060, 17616, 16960, 17066, 17034, 16113, 15246, 15743, 16570, 15383, 15784, 17132, 16029, 16049, 16903, 17405, 17475, 17765, 17661, 17717, 17680, 17716, 17660, 17860, 18320, 18572, 18097, 18032, 17589, 15921, 14980, 15054, 15033, 15140, 16526, 13353, 10618, 15439, 16819, 16681, 16398, 15656, 16736, 16983, 17792, 19086, 17095, 16842, 18838, 17748, 17796, 17886, 18139, 18496, 18178, 18269, 17407, 16940, 17342, 17239, 15912, 14954, 15222, 15109, 15136, 15184, 15029, 15598, 16415, 17089, 17636, 18048, 18791, 17820, 17721, 18177, 17058, 16788, 17769, 18406, 18055, 17898, 16939, 16416, 15497, 13603, 14502, 14278, 15185, 14619, 13733, 15205, 15537, 16479, 15931, 15313, 16704, 17438, 17835, 17097, 15877, 14594, 16431, 18264, 17037, 17322, 17181, 17167, 17351, 16930, 17808, 15045, 12894, 12793, 13546, 14110, 12176, 10790, 13836, 17425, 15847, 15136, 13414, 13862, 14867, 15067, 16260, 16048, 14548, 16361, 18112, 17303, 17213, 17507, 17628, 17411, 17414, 16276, 16212, 15062, 13954, 12458, 12290, 12812, 10822, 13126, 16335, 17302, 15525, 14296, 14607, 14526, 14441, 14723, 14086, 16224, 18269, 17334, 17375, 17076, 17724, 17604, 17275, 17266, 17348, 15843, 13985, 15081, 14478, 14844, 13655, 13911, 16738, 16893, 17977, 16885, 15335, 16273, 16740, 17285, 18492, 18491, 18002, 18105, 18475, 18117, 17811, 17633, 17935, 17581, 17696, 16669, 16406, 17296, 16970, 17139, 17051, 17086, 17081, 17209, 18090, 16558, 14379, 13579, 15512, 17210, 17202, 14957, 15364, 18369, 18080, 18562, 18350, 18228, 18611, 18019, 17835, 17374, 16867, 16650, 15941, 16107, 16678, 16272, 16083, 15410, 16690, 17332, 16519, 15884, 15363, 15054, 16548, 17279, 16660, 15713, 16437, 18564, 17841, 18216, 17994, 18153, 17990, 18223, 17192, 16175, 16085, 16095, 16032, 16423, 16627, 16036, 15876, 16265, 16877, 16682, 16139, 16147, 16167, 17701, 18223, 17249, 18594, 19373, 19811, 19952, 19605, 19665, 18873, 18260, 17844, 18564, 17596, 16249, 16597, 16242, 16554, 16483, 15998, 15924, 15965, 15802, 15844, 15857, 15783, 15947, 15608, 16681, 17591, 17964, 19396, 19880, 19763, 19132, 19458, 19256, 17883, 17782, 18291, 17106, 15893, 17079, 17446, 17765, 17078, 16026, 15909, 16355, 17300, 17428, 16956, 17340, 18382, 18010, 18212, 18405, 18846, 19310, 19805, 19449, 19257, 18809, 18539, 18562, 17917, 17967, 17933, 17914, 17995, 17824, 18173, 17054, 15949, 15693, 15648, 16941, 17157, 16957, 17892, 18463, 18091, 18349, 18712, 18970, 18792, 18313, 18964, 19168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 75, 0, 327, 0, 2770, 6270, 5629, 0, 10661, 24447, 17811, 19006, 19355, 19646, 19980, 20235, 20679, 21353, 21611, 21753, 21756, 21986, 22034, 22426, 22159, 21898, 22147, 21543, 22148, 22492, 24410, 26015, 25737, 25488, 26324, 24583, 28178, 16344, 4833, 8428, 6593, 6552, 7611, 8549, 4108, 632, 3266, 2319, 0, 324, 0, 91, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 166, 0, 576, 0, 8443, 8730, 7098, 22821, 26982, 26424, 26509, 26703, 26127, 27444, 22951, 18922, 21343, 20781, 21230, 21519, 22905, 23671, 23448, 23399, 23198, 22542, 22695, 22738, 25128, 27074, 25322, 25960, 23176, 24912, 12790, 3700, 8316, 7956, 8945, 4867, 5206, 5986, 5111, 3746, 3574, 1577, 0, 196, 0, 54, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 174, 0, 554, 0, 5199, 12994, 1916, 5313, 22010, 27454, 27960, 27468, 27463, 26800, 23059, 21250, 21225, 20984, 19712, 19163, 19173, 18763, 18107, 17169, 17859, 18692, 20813, 21527, 24366, 26665, 25340, 28365, 30588, 30068, 30126, 30475, 29568, 31511, 25536, 21279, 16147, 7399, 4923, 311, 75, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 294, 0, 1040, 0, 8931, 21965, 16425, 12226, 21437, 30903, 29576, 30227, 29736, 28170, 26731, 27242, 26845, 27329, 26553, 28018, 23431, 19770, 21580, 21012, 21954, 21957, 22336, 22771, 24640, 27616, 28873, 26922, 28504, 28949, 29880, 23396, 14565, 7326, 2179, 3496, 1657, 1788, 1404, 1757, 811, 0, 236, 266, 120, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 35, 0, 93, 765, 9327, 12286, 13119, 24147, 29733, 30656, 31220, 30030, 32372, 27234, 37030, 10691, 13284, 36475, 33755, 17856, 0, 4576, 122, 1833, 1801, 1645, 1730, 3958, 2798, 2471, 2253, 5341, 0, 18031, 31694, 23601, 25727, 22468, 23920, 23467, 23181, 24253, 22038, 26537, 11743, 0, 1458, 0, 417, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 216, 0, 778, 0, 5941, 12045, 11512, 15774, 18464, 26572, 30758, 31092, 31141, 31175, 30307, 29069, 26263, 24898, 24061, 22585, 22786, 22689, 22605, 22975, 22125, 23882, 22341, 33055, 17070, 0, 4778, 1280, 4412, 1885, 5695, 0, 16400, 34338, 21858, 22097, 19843, 21733, 9119, 0, 1501, 0, 328, 0, 3008, 5137, 5295, 5962, 6283, 6140, 6914, 2769, 0, 322, 0, 59, 268, 2222, 3583, 3399, 3354, 3273, 3442, 3125, 3762, 1666, 0, 206, 0, 59, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 353, 0, 1275, 0, 9351, 17532, 18463, 30582, 30982, 31375, 27701, 24183, 20862, 19427, 20510, 19734, 19898, 20062, 21080, 21131, 22754, 25385, 26120, 26485, 26731, 28236, 27219, 29519, 28584, 36394, 15409, 201, 545, 17031, 32934, 26218, 30123, 23444, 23860, 21479, 18098, 6727, 657, 2318, 1469, 1997, 1594, 2053, 876, 0, 111, 0, 31, 0, 1, 5, 0, 41, 0, 144, 0, 1311, 4248, 4409, 4212, 2587, 8190, 4959, 0, 678, 0, 194, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 173, 0, 558, 0, 4903, 13632, 10760, 12193, 4752, 14757, 26826, 24124, 22492, 17886, 20167, 19542, 19687, 19751, 19643, 19596, 19744, 19678, 19460, 19679, 21084, 21918, 21980, 22161, 22032, 22210, 21909, 22467, 21345, 24946, 28216, 29992, 30717, 32290, 24487, 20713, 13511, 2448, 2781, 6145, 10501, 8753, 5454, 2112, 4543, 5401, 5458, 5418, 4968, 5741, 2480, 0, 305, 0, 83, 0, 0, 34, 0, 152, 0, 1194, 2653, 2411, 1643, 111, 23, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 336, 0, 1172, 0, 9465, 21532, 17930, 20160, 19409, 20137, 19972, 20464, 21598, 22190, 22062, 22117, 22121, 20881, 21115, 22280, 21191, 24536, 27609, 25388, 26336, 24396, 26775, 11514, 0, 5821, 5471, 7860, 4281, 4915, 6558, 5395, 5509, 5299, 6497, 1318, 2152, 5535, 3738, 4605, 4057, 4504, 3985, 4852, 2140, 0, 266, 0, 76, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 301, 0, 1097, 0, 7512, 10349, 7680, 17157, 20731, 20823, 17866, 19375, 18926, 18983, 18990, 18337, 17932, 18150, 18433, 20121, 22128, 20898, 21649, 21947, 20112, 20713, 19240, 22693, 25420, 24179, 24780, 24368, 24768, 24213, 25221, 22422, 20291, 12323, 10417, 16117, 16797, 6793, 0, 808, 0, 222, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 266, 0, 901, 0, 7292, 16404, 10411, 9532, 3061, 0, 333, 0, 100, 0, 1, 12, 0, 579, 3188, 3345, 3013, 4316, 6446, 9381, 2366, 2476, 10166, 6420, 1123, 46, 1847, 3623, 4741, 4817, 4994, 3087, 1195, 1408, 399, 0, 34, 0, 11, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 139, 0, 578, 0, 4213, 6953, 7073, 0, 10925, 29291, 27497, 30505, 29671, 29981, 29018, 29269, 28813, 29797, 27399, 35940, 16655, 0, 3612, 938, 3863, 2983, 4082, 3826, 3819, 3908, 3381, 4735, 4832, 3975, 4826, 5298, 4278, 3793, 3937, 3715, 4123, 3374, 4773, 1939, 11412, 21981, 21526, 21747, 24236, 11863, 343, 3829, 2984, 5373, 4990, 5905, 2233, 0, 213, 0, 0, 283, 0, 2525, 5830, 5616, 11457, 5155, 0, 632, 0, 190, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 142, 0, 1656, 951, 10110, 19968, 18014, 15332, 23704, 31568, 27623, 26932, 21899, 18646, 19994, 20518, 21417, 21528, 21757, 21255, 22268, 20146, 27157, 33304, 30704, 26523, 33761, 16065, 0, 6029, 3735, 6255, 3701, 6974, 0, 16898, 32178, 22989, 24782, 21653, 21318, 18871, 17965, 14925, 8906, 6678, 6643, 4879, 1576, 0, 165, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 220, 0, 745, 0, 6599, 18317, 17606, 17449, 11782, 9501, 14771, 18037, 19353, 19555, 21088, 22368, 22564, 22925, 22693, 24015, 25719, 26164, 26197, 26496, 26675, 25367, 23683, 23390, 22487, 24233, 24640, 26125, 25856, 31745, 14293, 0, 6574, 5039, 5609, 5498, 5927, 5360, 4792, 5041, 4818, 5118, 4621, 5580, 2466, 0, 306, 0, 87, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 201, 0, 739, 0, 6289, 7752, 10043, 25571, 29380, 27964, 25182, 23136, 22001, 22963, 23318, 25077, 28278, 30227, 28998, 28219, 29508, 30867, 31478, 31423, 31230, 31723, 30743, 32735, 26568, 23168, 26307, 25041, 26694, 32204, 23471, 8070, 6915, 7042, 6264, 4719, 2746, 1283, 1628, 1246, 387, 0, 38, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 303, 0, 1058, 0, 8665, 20427, 18094, 20105, 19299, 19518, 19531, 20414, 20859, 23993, 24168, 22039, 22384, 22058, 22078, 21939, 22915, 23723, 24363, 23347, 25561, 23895, 25455, 10384, 0, 1804, 11496, 25290, 21153, 24882, 12387, 4633, 5088, 548, 2366, 454, 0, 23, 0, 19, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 71, 0, 127, 0, 3120, 14620, 3123, 8736, 27861, 26540, 26940, 20617, 19423, 20666, 20358, 20788, 20514, 20586, 20632, 21010, 21447, 21598, 21847, 21762, 21614, 21712, 21684, 21135, 20056, 19449, 19770, 19304, 20149, 18562, 21759, 11908, 4748, 4570, 15122, 15759, 4210, 6259, 3188, 4389, 2948, 1357, 54, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 34, 0, 120, 0, 791, 791, 0, 120, 0, 34, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 156, 0, 441, 0, 4605, 13047, 416, 9381, 23311, 19751, 21691, 20611, 21200, 20879, 21086, 20781, 20851, 21069, 21268, 21521, 21502, 21463, 21414, 20808, 19842, 19758, 19531, 19245, 19774, 20196, 22417, 26060, 9373, 0, 2470, 4564, 5722, 6112, 6245, 3193, 2828, 3567, 2308, 1844, 2317, 438, 0, 17, 0, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 140, 0, 542, 0, 4467, 10177, 9820, 5704, 16159, 26542, 22104, 21286, 19370, 20456, 20122, 20834, 20865, 21868, 22682, 22687, 22418, 21763, 21901, 21942, 21823, 21634, 20678, 19560, 19803, 19547, 20109, 20072, 24002, 25830, 26170, 29641, 29740, 30008, 29619, 30295, 29047, 31468, 24898, 24278, 17019, 5217, 9596, 6269, 1721, 0, 144, 0, 27, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 208, 0, 726, 0, 5144, 7295, 0, 428, 0, 449, 0, 1211, 0, 9764, 22779, 19920, 21993, 21525, 22500, 22355, 22727, 22712, 22649, 22462, 22175, 22245, 23415, 24310, 23310, 25596, 26765, 26232, 25788, 23704, 16963, 7635, 6302, 7609, 7176, 6710, 6406, 7174, 5756, 7187, 2159, 2006, 3172, 0, 534, 0, 141, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 67, 0, 367, 0, 2527, 4719, 13051, 4192, 10784, 29093, 24098, 26087, 20160, 17323, 17202, 16831, 18728, 18935, 19739, 20509, 20471, 21245, 20590, 21306, 21444, 21458, 22101, 22409, 23052, 23038, 24725, 25449, 25467, 25105, 25918, 24354, 27546, 16493, 2581, 6881, 5338, 4850, 6118, 4775, 3875, 3289, 3763, 1595, 0, 195, 0, 55, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 177, 0, 626, 0, 5133, 11085, 6938, 10189, 20974, 26192, 24857, 25469, 25169, 25283, 25329, 24758, 22907, 21717, 21796, 21622, 20769, 19538, 18524, 17945, 17132, 18053, 17520, 21334, 23863, 25448, 23968, 28939, 16337, 0, 17037, 29176, 18510, 20774, 21296, 20770, 17421, 8941, 3959, 2282, 166, 27, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 86, 0, 295, 0, 3131, 3702, 137, 346, 0, 79, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 285, 0, 1000, 0, 8638, 21538, 16159, 13261, 21636, 29575, 27952, 27925, 26789, 25580, 23915, 23225, 23805, 24172, 23845, 24263, 24481, 22682, 21847, 22376, 21432, 21471, 22574, 22382, 23591, 23228, 26782, 29437, 27664, 27730, 28779, 30304, 30046, 30513, 29690, 31192, 28428, 33954, 15838, 0, 3759, 3016, 1805, 539, 1535, 0, 247, 0, 65, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 253, 0, 945, 0, 6519, 10420, 13944, 25681, 28057, 32194, 31111, 30982, 31465, 30255, 29709, 29825, 30064, 29389, 30761, 28172, 33372, 16262, 0, 4464, 2037, 3327, 1018, 283, 1589, 3123, 2313, 5910, 0, 15922, 28910, 21228, 24678, 21842, 20743, 17218, 15885, 5692, 0, 1890, 283, 9, 0, 0, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 233, 0, 832, 0, 8584, 15103, 13898, 16241, 15719, 26192, 30702, 30147, 30385, 29296, 28610, 24131, 21064, 22914, 23700, 24064, 24287, 25235, 25568, 26515, 27110, 26742, 22008, 30960, 14769, 0, 4459, 2351, 3381, 3214, 2311, 5740, 0, 16484, 33165, 20601, 21438, 19858, 20597, 19805, 20928, 18981, 22838, 10127, 0, 1327, 0, 609, 0, 2378, 5308, 4453, 1633, 0, 191, 0, 43, 0, 0, 46, 0, 431, 916, 205, 0, 11, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 109, 0, 285, 0, 6813, 14298, 2704, 6514, 16818, 24501, 28628, 25815, 22844, 18460, 20331, 19622, 20177, 20028, 20077, 19546, 20887, 22736, 22753, 22866, 22753, 22907, 22645, 23405, 24383, 26457, 29972, 21105, 5804, 0, 8703, 20494, 17892, 24042, 25245, 19309, 21316, 9423, 73, 2624, 1142, 1863, 1111, 1456, 668, 2039, 1424, 0, 203, 0, 57, 0, 8, 0, 0, 12, 0, 40, 0, 529, 2310, 2902, 2807, 2791, 2903, 2651, 3183, 1411, 0, 175, 0, 50, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 444, 0, 1528, 0, 12570, 29134, 21075, 21415, 20551, 20206, 20400, 20804, 21911, 22864, 22010, 20933, 20173, 20059, 21233, 21651, 22336, 22609, 23121, 22749, 22388, 22728, 26561, 27107, 29304, 24449, 36625, 11837, 12431, 32358, 18405, 15362, 683, 9547, 7855, 3459, 4908, 3653, 3751, 3655, 3626, 3799, 3442, 4155, 1836, 0, 228, 0, 65, 0, 15, 0, 3, 0, 5, 0, 215, 1215, 629, 0, 79, 0, 23, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 169, 0, 609, 0, 5043, 11506, 8686, 9353, 18424, 25092, 20603, 19614, 20746, 20246, 19514, 19842, 20585, 20759, 21399, 21606, 21527, 22525, 23007, 22724, 22561, 22456, 22291, 22326, 22314, 22354, 22236, 22410, 23382, 29925, 13897, 584, 7040, 7111, 6142, 5435, 6679, 5612, 5473, 5626, 5895, 2697, 0, 3110, 2710, 0, 394, 0, 114, 0, 23, 0, 0, 0, 12, 0, 70, 0, 251, 0, 1636, 1768, 504, 1498, 148, 23, 0, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 108, 0, 402, 0, 3263, 8287, 10921, 9534, 6251, 7205, 6987, 6627, 7691, 5334, 13221, 20697, 17091, 17659, 17872, 18035, 18690, 20588, 21601, 22497, 22831, 22892, 22770, 21396, 24754, 27469, 26540, 26170, 25993, 27972, 27355, 28766, 22716, 18932, 18591, 16769, 10491, 2246, 9827, 17831, 6687, 0, 722, 0, 212, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 194, 0, 652, 0, 5627, 14169, 10684, 15431, 20151, 26367, 31605, 31006, 29323, 26233, 25747, 25253, 24053, 21830, 20001, 19160, 17990, 17059, 16860, 17005, 17730, 20941, 20439, 20182, 21522, 23296, 9112, 0, 1192, 0, 402, 113, 7, 836, 763, 0, 114, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 69, 0, 246, 0, 2371, 6117, 3086, 5315, 20523, 29512, 28601, 28644, 28370, 28769, 28794, 28743, 29059, 28334, 29728, 27135, 32319, 15339, 0, 4410, 2687, 4694, 3774, 4118, 4432, 4055, 4762, 5849, 5067, 4224, 4450, 5807, 2915, 5979, 0, 16849, 28077, 13592, 12872, 11895, 20924, 21528, 22641, 22497, 24155, 12068, 1363, 4509, 2081, 2996, 1196, 0, 149, 0, 49, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 107, 0, 919, 2625, 4899, 6479, 11027, 15231, 10757, 16384, 17393, 22640, 32650, 31597, 29999, 26910, 28129, 29184, 27051, 29538, 28389, 35848, 16677, 0, 2945, 270, 2264, 1849, 1462, 407, 1449, 3044, 5192, 5580, 6206, 4413, 6772, 0, 17345, 31507, 20871, 23916, 21883, 23331, 21930, 24025, 17697, 10649, 8591, 5628, 2663, 0, 343, 0, 68, 0, 11, 0, 0, 2, 0, 7, 0, 48, 48, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 48, 804, 9684, 17132, 14771, 12681, 12771, 17938, 19731, 19390, 20965, 20918, 22283, 23279, 22395, 22876, 24569, 24889, 25048, 24984, 25024, 24979, 25066, 24825, 24789, 23722, 25860, 25196, 28073, 25582, 28123, 22475, 4738, 6023, 6671, 5903, 5880, 5371, 6253, 2786, 0, 276, 0, 80, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 91, 0, 311, 0, 4518, 21651, 29986, 27232, 26287, 23426, 21601, 22474, 23258, 24759, 26650, 29201, 28551, 28183, 28551, 29274, 30618, 32194, 28870, 24254, 23381, 22823, 22908, 23958, 24346, 25773, 26804, 26395, 28795, 33680, 26341, 10955, 7256, 6709, 4229, 2396, 1626, 1422, 1405, 1423, 1393, 1463, 1329, 1601, 708, 0, 88, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 79, 0, 193, 0, 2924, 14305, 14056, 14012, 2957, 8019, 23883, 18971, 20401, 19822, 20120, 20267, 20059, 20218, 20811, 23727, 26347, 26377, 25262, 23965, 24027, 24174, 24087, 24217, 23997, 24347, 23724, 25495, 22633, 6170, 799, 3523, 13745, 24682, 16423, 6988, 4821, 3060, 1240, 1833, 630, 0, 57, 0, 20, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 0, 60, 0, 413, 773, 1408, 826, 0, 113, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 227, 0, 795, 0, 6275, 13471, 10596, 11832, 11356, 11262, 11958, 10276, 15980, 21507, 19759, 20802, 21016, 21713, 21624, 22592, 23379, 23601, 23739, 22742, 22865, 22989, 22303, 22693, 21962, 22145, 21276, 23456, 25652, 27495, 15101, 5703, 9570, 7052, 6936, 7094, 6448, 5308, 4753, 4200, 3671, 1571, 54, 26, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 21, 0, 76, 0, 503, 503, 0, 76, 0, 21, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 157, 0, 448, 0, 4699, 13419, 716, 9243, 24830, 22401, 21476, 18851, 20266, 20151, 20048, 19616, 20129, 21983, 22394, 22076, 22625, 22831, 22464, 22018, 22242, 21769, 21172, 21287, 21222, 21467, 21834, 21887, 22047, 21666, 22409, 21025, 23809, 14420, 3114, 3945, 1652, 1924, 1048, 1937, 2709, 730, 0, 60, 0, 20, 0, 5, 0, 0, 0, 0, 8, 0, 49, 0, 179, 0, 2482, 6059, 7751, 8517, 7963, 5759, 1133, 0, 74, 0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 0, 88, 0, 1656, 8902, 14112, 1047, 9360, 25781, 19403, 19148, 20036, 20332, 20259, 20315, 20199, 20451, 19900, 21727, 23545, 23047, 23339, 23535, 23585, 23510, 23609, 22828, 22595, 22597, 22585, 23567, 26831, 28001, 29582, 25642, 21217, 10095, 938, 6448, 7049, 7592, 11526, 16920, 17785, 16577, 20966, 10799, 0, 540, 0, 169, 0, 29, 0, 0, 0, 17, 0, 85, 0, 301, 0, 2340, 4790, 3198, 1306, 0, 167, 0, 42, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29729, 28756, 29021, 29343, 30109, 29864, 29423, 27373, 27753, 17661, 9426, 11332, 9064, 6439, 4361, 4827, 3119, 6387, 7639, 6223, 6971, 6350, 6710, 6393, 6799, 6141, 7409, 3277, 0, 407, 0, 116, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 154, 0, 533, 0, 4646, 12324, 11273, 11319, 11286, 11074, 11622, 10547, 12711, 5620, 0, 698, 0, 199, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 199, 200, 0, 32, 0, 0, 120, 0, 460, 0, 1583, 0, 12871, 29604, 30924, 29377, 37992, 12439, 11661, 38288, 26198, 29305, 27240, 27839, 26824, 27092, 27547, 27691, 27848, 27791, 27466, 26958, 27007, 27175, 27125, 26867, 27139, 27334, 27275, 27427, 27171, 27349, 27232, 27054, 27219, 27327, 27337, 27250, 27077, 26895, 26884, 26871, 26897, 26849, 26936, 26761, 27369, 28269, 28450, 28514, 28168, 28312, 28849, 28833, 28558, 27444, 25123, 9013, 0, 718, 0, 164, 0, 0, 264, 0, 3131, 8342, 8559, 11200, 6975, 5279, 3148, 0, 458, 0, 123, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 449, 634, 1453, 3341, 8059, 11616, 11241, 12403, 12264, 12519, 13705, 12100, 9592, 8656, 8837, 8839, 8689, 9062, 8007, 8427, 9288, 9248, 6665, 1094, 0, 43, 0, 17, 0, 10, 0, 17, 0, 182, 572, 215, 0, 42, 0, 102, 0, 348, 0, 2802, 6309, 5676, 5441, 8896, 17607, 22605, 24389, 24662, 24549, 24327, 24527, 24536, 24866, 25144, 25219, 24849, 25715, 23906, 28525, 28250, 34547, 17061, 0, 4842, 0, 15828, 33760, 28054, 29080, 26896, 29104, 28852, 29727, 29780, 30184, 29896, 29055, 28604, 27906, 26215, 25357, 24622, 24492, 22413, 20564, 20555, 20388, 21069, 22742, 23853, 23174, 22578, 21262, 18240, 15194, 5986, 317, 1920, 1104, 1598, 1240, 1620, 688, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 97, 0, 788, 1770, 1488, 1597, 1597, 1488, 1770, 763, 0, 0, 180, 0, 815, 0, 7184, 19632, 23131, 28363, 30291, 31653, 31480, 31327, 31073, 30188, 28701, 28755, 29537, 30297, 29666, 24109, 6843, 0, 652, 0, 126, 0, 0, 387, 0, 3492, 10080, 17192, 25593, 26916, 28239, 28799, 28649, 28748, 28657, 28757, 28596, 29041, 29288, 29100, 29251, 28884, 29315, 27386, 30344, 24922, 36642, 12715, 11229, 35291, 26052, 25004, 17195, 20176, 18045, 17535, 17110, 16819, 16744, 15639, 13810, 13981, 12987, 12027, 11634, 13314, 17201, 20289, 18056, 10091, 0, 21398, 20210, 0, 3028, 0, 862, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 98, 0, 860, 3663, 12413, 19618, 21657, 23747, 25181, 29501, 26490, 34020, 15395, 0, 3124, 474, 2480, 1666, 2125, 2079, 1655, 2143, 177, 2689, 0, 14922, 33484, 27753, 30665, 28562, 28927, 28694, 28846, 28728, 29147, 29912, 29825, 29906, 29877, 30477, 30977, 30853, 30866, 30947, 30742, 31186, 29700, 28311, 29043, 28972, 28897, 29420, 28322, 27350, 27860, 27950, 28367, 28566, 28565, 29118, 29502, 29510, 29114, 26687, 25628, 23871, 22411, 18998, 15932, 17227, 13943, 3746, 0, 365, 0, 206, 0, 1000, 2973, 5729, 6937, 8708, 6826, 4477, 5936, 5318, 5624, 5492, 5502, 5634, 4718, 1237, 0, 110, 0, 32, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 63, 0, 217, 0, 3282, 16384, 24411, 26399, 27429, 27619, 28452, 28576, 28789, 28482, 29244, 28456, 30417, 26234, 35154, 11226, 11131, 35139, 26550, 30665, 27823, 28655, 28226, 28069, 28043, 27924, 27671, 27087, 26727, 26555, 25993, 25995, 25918, 25756, 25848, 25735, 25911, 25583, 26667, 27935, 27699, 28624, 28757, 29185, 29460, 29372, 29122, 28990, 29295, 29199, 29462, 28562, 28209, 28308, 28284, 28496, 27945, 26225, 25554, 25371, 24331, 19696, 19266, 7730, 0, 935, 0, 311, 0, 219, 0, 1337, 2965, 2562, 3140, 3477, 3217, 2823, 2880, 2964, 2720, 3257, 1446, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 181, 0, 644, 0, 5590, 15414, 18416, 21927, 22115, 23000, 24139, 24678, 26925, 28990, 29354, 30287, 30529, 31270, 32736, 30316, 28103, 28985, 28669, 28927, 28812, 28898, 29066, 29242, 29244, 29119, 29017, 29002, 29109, 29060, 29175, 29091, 29070, 29080, 29416, 29604, 29615, 29759, 29691, 29741, 29677, 29798, 29551, 30079, 28237, 22424, 6732, 0, 688, 0, 195, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 105, 0, 370, 0, 2940, 6755, 6916, 9300, 8598, 10484, 11568, 10073, 10178, 8487, 6650, 7166, 4528, 2479, 3100, 2730, 3041, 2677, 3275, 1438, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 294, 0, 1019, 0, 8470, 19456, 15891, 19699, 27043, 26961, 34882, 17080, 0, 4858, 0, 16487, 33604, 27260, 30332, 28353, 29267, 28868, 29213, 29250, 29259, 29179, 28921, 29078, 29193, 29152, 29192, 29134, 29232, 29046, 29598, 29849, 29653, 29836, 29886, 29789, 29651, 30125, 29869, 29617, 28734, 27427, 24015, 25256, 14999, 773, 261, 0, 92, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 86, 0, 310, 0, 2330, 4340, 3446, 3700, 3914, 1910, 0, 246, 0, 66, 0, 0, 63, 0, 353, 0, 1250, 0, 9978, 22754, 22543, 27475, 26185, 26737, 26772, 27588, 27786, 27843, 27737, 27664, 27731, 28081, 28284, 28306, 27896, 27048, 26932, 25972, 25259, 25477, 25342, 25465, 25298, 25601, 24666, 23170, 20579, 22430, 26477, 27644, 28501, 28471, 28440, 28706, 28207, 29436, 26860, 32802, 14354, 0, 3843, 1917, 2013, 4528, 0, 16727, 36685, 30362, 32253, 29576, 30273, 29576, 28382, 23000, 19920, 17664, 12005, 10252, 10627, 10158, 9609, 9073, 9185, 8922, 9402, 8527, 10275, 4546, 0, 564, 0, 161, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 134, 0, 521, 0, 7059, 23692, 28677, 30816, 29245, 36487, 16512, 0, 4430, 1399, 3171, 2226, 2136, 1707, 1881, 1879, 2312, 2663, 2873, 2916, 3086, 3002, 3038, 3088, 2942, 2827, 2961, 3092, 2779, 2965, 2902, 3214, 4256, 4613, 4466, 4717, 4184, 5250, 3232, 7135, 0, 14695, 32988, 26711, 30097, 28528, 29147, 28531, 28844, 29161, 29286, 28761, 30004, 28750, 28815, 19800, 3371, 0, 149, 0, 47, 0, 5, 0, 0, 68, 0, 239, 0, 2139, 6099, 7060, 7983, 8212, 8006, 8398, 8053, 7153, 7533, 7188, 7647, 6899, 8333, 3683, 0, 457, 0, 130, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2607, 2603, 2628, 2569, 2733, 2595, 2206, 2342, 2401, 1956, 1903, 2367, 2721, 2677, 2807, 2675, 2664, 1122, 0, 264, 0, 1111, 2469, 2648, 2983, 3133, 1637, 0, 1595, 1326, 0, 191, 0, 59, 0, 27, 0, 52, 0, 462, 1199, 809, 613, 705, 575, 799, 362, 1792, 3362, 3154, 3294, 2794, 2730, 2959, 2728, 3167, 3662, 3459, 3569, 3536, 3573, 3634, 3644, 3658, 3579, 3514, 3486, 3554, 3510, 3727, 3335, 3145, 1245, 0, 149, 0, 42, 0, 8, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1285, 2965, 2562, 2868, 2825, 3209, 3370, 3459, 3301, 3306, 2863, 2350, 2397, 2337, 2322, 2327, 2576, 2591, 2584, 2690, 2645, 3075, 3563, 3646, 3751, 3739, 3663, 3749, 3920, 3879, 3913, 4017, 3943, 3919, 3406, 3743, 1539, 0, 185, 0, 57, 0, 33, 0, 77, 0, 699, 2015, 2095, 2642, 2848, 2892, 2953, 3145, 3297, 3609, 3911, 3813, 3824, 3669, 3908, 3479, 2772, 2703, 2764, 2793, 2432, 3042, 3115, 2604, 2838, 2847, 3127, 2943, 3608, 4324, 3625, 3641, 3807, 3733, 3743, 3834, 3976, 3925, 3959, 3927, 3967, 3907, 4008, 3547, 2777, 3064, 994, 0, 0, 1423, 3447, 2926, 3416, 3358, 3478, 3283, 3430, 3599, 3668, 3843, 3766, 3720, 3149, 2812, 2975, 2935, 2870, 2950, 2861, 2872, 3102, 3003, 2992, 2901, 2927, 2895, 2841, 2861, 2850, 2955, 2962, 2955, 2976, 2933, 3015, 2850, 3389, 3918, 3746, 3861, 3996, 3990, 3979, 3832, 3529, 3766, 3722, 3507, 3274, 3164, 3274, 3391, 3493, 3466, 3450, 3387, 3551, 3630, 3747, 3890, 4122, 3965, 3821, 3441, 2928, 2930, 2705, 2616, 2702, 2742, 2715, 2850, 2728, 2730, 2849, 2807, 2829, 2818, 2822, 2823, 2826, 2891, 2891, 3252, 3685, 3601, 3812, 4042, 3996, 4113, 4198, 4253, 4290, 4082, 4147, 4156, 3827, 4136, 3845, 3307, 3282, 3287, 3437, 3434, 3410, 3289, 3320, 3279, 3532, 3670, 3673, 3894, 3721, 3713, 3101, 2719, 2902, 2689, 2656, 2650, 2661, 2643, 2677, 2608, 2838, 3095, 3111, 3125, 2975, 2869, 2700, 2676, 2797, 2596, 2995, 3471, 3481, 3466, 3472, 3755, 3746, 4134, 4552, 4617, 4603, 4528, 4531, 4538, 4169, 3749, 3590, 3277, 3268, 3285, 3134, 3157, 3377, 3340, 3264, 3413, 3301, 3450, 3619, 3576, 3581, 3610, 3536, 3695, 3165, 2649, 2928, 2952, 3180, 3119, 3111, 3174, 2888, 2862, 2932, 2823, 2864, 2804, 3206, 3626, 3560, 3600, 3713, 3672, 3748, 3837, 4291, 4683, 4653, 4774, 4883, 4740, 4700, 4885, 5380, 2045, 0, 290, 0, 756, 2622, 2718, 2278, 2407, 2365, 2350, 2431, 2234, 2895, 3500, 3467, 3446, 3447, 3647, 3593, 3175, 2997, 3301, 3184, 3157, 3320, 3198, 2691, 2536, 2610, 2418, 2361, 2750, 2747, 3149, 3461, 3451, 3564, 3548, 3800, 4020, 4158, 4504, 4849, 4687, 4894, 4166, 3446, 3532, 3541, 3850, 3828, 3897, 3775, 3999, 3583, 4412, 1830, 41, 598, 0, 0, 947, 2332, 1968, 2535, 2698, 2807, 2958, 3171, 3322, 3199, 3096, 3198, 2794, 2611, 2813, 2776, 2347, 1898, 1901, 2134, 2126, 2084, 2933, 2866, 2888, 3471, 3461, 3613, 3825, 4131, 4195, 4327, 3985, 3692, 3772, 3744, 3738, 3781, 3682, 4025, 4386, 3910, 4106, 3937, 4670, 1999, 0, 239, 0, 361, 808, 205, 482, 1898, 1875, 2311, 2894, 2946, 3043, 3215, 3393, 3523, 3572, 3459, 3339, 2995, 3055, 1274, 0, 767, 1422, 1478, 1894, 2663, 3082, 3007, 3337, 3503, 3459, 3485, 3461, 3492, 3440, 3573, 3593, 3728, 4011, 4047, 4270, 4041, 3832, 4474, 4037, 4667, 2051, 0, 255, 0, 73, 0, 14, 0, 3, 0, 13, 0, 219, 1263, 2507, 2984, 3053, 3159, 3215, 3334, 3269, 3369, 3078, 2862, 1212, 0, 907, 1695, 1482, 1623, 1477, 1681, 1317, 2487, 3844, 3758, 3918, 3700, 3683, 3446, 3580, 3842, 3840, 3897, 4077, 3828, 3718, 4283, 4141, 4540, 1782, 0, 210, 0, 60, 0, 11, 0, 0, 7, 0, 30, 0, 239, 707, 1827, 2918, 3003, 3113, 3176, 3358, 3414, 3410, 3395, 3432, 3355, 3514, 2998, 2459, 2374, 2762, 3302, 3082, 3322, 3634, 3645, 3789, 3856, 3449, 3671, 3451, 3731, 4101, 3861, 4196, 4136, 4151, 4298, 3821, 3647, 1364, 0, 158, 0, 45, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 57, 0, 198, 0, 1686, 4066, 2623, 1909, 2272, 1094, 0, 958, 2602, 805, 467, 2357, 2648, 2860, 3129, 3519, 3621, 3925, 3868, 3623, 1226, 0, 134, 0, 38, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 43, 0, 151, 0, 1261, 3067, 2818, 3081, 3277, 3727, 3720, 3753, 3682, 3550, 2851, 2622, 3014, 2730, 2714, 2732, 2528, 1975, 1991, 2294, 2362, 2488, 2958, 3456, 3499, 3642, 3758, 3739, 3526, 1189, 0, 129, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1309, 3083, 2367, 2857, 3328, 3503, 3485, 3527, 3674, 2519, 2170, 2806, 2438, 2502, 2931, 2804, 2836, 2952, 2985, 2783, 2548, 2848, 2134, 2085, 2400, 2392, 2706, 2688, 3101, 3333, 3467, 3700, 3724, 3817, 3699, 3902, 3536, 4262, 1885, 0, 234, 0, 62, 0, 0, 38, 0, 157, 0, 1291, 3082, 2892, 3351, 3233, 3409, 3391, 3439, 3183, 2353, 2047, 2147, 2106, 2471, 2617, 2601, 2867, 2904, 2945, 2904, 2999, 2993, 3037, 3100, 3113, 3177, 3157, 3190, 3172, 3191, 3163, 3217, 3105, 3458, 3711, 3875, 3631, 4087, 1743, 0, 213, 0, 60, 0, 23, 0, 55, 0, 198, 0, 1535, 3184, 2688, 3264, 3338, 3279, 3075, 3388, 3417, 806, 746, 2671, 2388, 2739, 2891, 3131, 3090, 3141, 3205, 3202, 3278, 3305, 3300, 3291, 3317, 3263, 3372, 3062, 2957, 2587, 2304, 2554, 2654, 2655, 3131, 3661, 3410, 3606, 3396, 3877, 1569, 0, 187, 0, 60, 0, 42, 0, 112, 0, 928, 2347, 2663, 3253, 3125, 3577, 3298, 3287, 3174, 2680, 2426, 2160, 2705, 2798, 2667, 2680, 2664, 2679, 2664, 2684, 2646, 2802, 3136, 2995, 2962, 3050, 3042, 3091, 2938, 2810, 2708, 2718, 2749, 2786, 2771, 2844, 2873, 3252, 3614, 3516, 3579, 3429, 3444, 2867, 2792, 1143, 0, 112, 0, 0, 155, 0, 1446, 3469, 3085, 3451, 3339, 3584, 3369, 3097, 3229, 3077, 3308, 2915, 3660, 1402, 435, 2659, 369, 867, 2333, 1965, 2349, 2473, 2462, 2161, 1735, 2102, 883, 0, 66, 15, 0, 698, 2162, 2158, 2713, 3194, 3264, 3542, 3490, 3727, 3390, 2665, 894, 0, 99, 0, 27, 0, 5, 0, 0, 9, 0, 39, 0, 120, 0, 1186, 3394, 1121, 0, 0, 445, 1575, 1813, 2313, 2622, 2539, 2648, 2853, 2764, 2505, 2510, 2230, 2159, 868, 0, 93, 0, 0, 276, 1447, 1971, 2544, 3068, 3161, 3364, 3536, 3491, 3645, 3341, 4500, 2102, 0, 265, 0, 76, 0, 12, 0, 0, 18, 0, 65, 0, 656, 2240, 2733, 2464, 2465, 2800, 2468, 2351, 768, 0, 0, 742, 2480, 2472, 2438, 2234, 2817, 1208, 0, 153, 0, 66, 0, 92, 0, 725, 1943, 2097, 2604, 3124, 3496, 3423, 3426, 3580, 3619, 3653, 3560, 3745, 3398, 4093, 1811, 0, 225, 0, 64, 0, 10, 0, 0, 35, 0, 133, 0, 857, 967, 1037, 2248, 2152, 2532, 2135, 2653, 1100, 0, 90, 10, 0, 536, 564, 0, 76, 0, 0, 34, 0, 405, 1063, 901, 1713, 2244, 2092, 2178, 2112, 2181, 2077, 2454, 3322, 3426, 3569, 3555, 4068, 1647, 0, 196, 0, 56, 0, 11, 0, 0, 0, 0, 0, 0, 0, 3, 0, 8, 0, 15, 0, 424, 2216, 1116, 0, 140, 0, 41, 0, 9, 0, 0, 0, 10, 0, 47, 0, 160, 0, 1413, 3532, 2204, 2589, 4061, 3174, 3091, 3816, 3322, 3472, 3740, 3682, 3620, 2885, 3672, 1737, 0, 221, 0, 63, 0, 12, 0, 0, 0, 3, 0, 13, 0, 46, 0, 427, 1188, 1080, 1652, 2702, 2678, 2118, 2012, 2045, 1989, 2092, 1903, 2278, 1029, 0, 187, 0, 673, 2148, 2633, 2571, 3284, 1190, 0, 0, 1661, 3948, 3076, 3473, 3550, 3427, 3819, 1552, 0, 184, 0, 53, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 93, 0, 787, 2019, 1704, 2587, 1112, 0, 79, 31, 0, 1002, 3045, 2246, 1954, 821, 0, 104, 0, 30, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 0, 42, 0, 554, 2079, 890, 0, 103, 0, 31, 0, 7, 0, 0, 6, 0, 24, 0, 74, 0, 778, 2400, 889, 0, 94, 0, 29, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 55, 0, 895, 1603, 389, 0, 27, 0, 9, 0, 3, 0, 0, 0, 0, 0, 2, 0, 5, 0, 12, 0, 288, 1449, 718, 0, 89, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 25, 0, 90, 0, 595, 595, 0, 90, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 198, 198, 0, 30, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 19, 0, 68, 0, 450, 450, 0, 68, 0, 19, 0, 3, 0, 0, 0, 0, 0, 1, 0, 5, 0, 19, 0, 125, 125, 0, 19, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 633, 1429, 2018, 2193, 2176, 2138, 2240, 2037, 2451, 1085, 0, 134, 0, 38, 0, 7, 0, 1, 0, 8, 0, 28, 0, 424, 321, 0, 46, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 44, 0, 147, 0, 1224, 2670, 631, 0, 40, 0, 15, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 47, 0, 175, 0, 1129, 962, 39, 1004, 2360, 3010, 2596, 2805, 692, 0, 56, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 60, 0, 218, 0, 1457, 1475, 0, 599, 1961, 1133, 0, 147, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 56, 0, 206, 0, 1345, 1250, 0, 0, 651, 815, 0, 126, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1545, 1610, 1540, 1582, 1739, 1395, 2115, 740, 3287, 0, 14847, 31206, 25333, 28322, 26995, 26416, 27153, 24572, 24692, 10264, 0, 1048, 0, 301, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 86, 338, 214, 277, 251, 66, 132, 97, 117, 104, 115, 85, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 883, 0, 3138, 0, 20590, 20829, 0, 4379, 0, 2528, 1622, 2417, 2410, 2739, 3011, 3195, 2770, 2929, 3393, 3468, 3258, 3103, 3078, 2897, 2915, 2764, 2726, 2823, 2505, 2027, 1547, 1459, 1358, 1269, 1416, 1452, 1526, 1480, 1541, 1439, 1621, 1260, 2459, 3790, 3566, 3594, 3562, 3830, 3453, 3247, 3190, 3149, 3104, 2694, 2150, 634, 0, 64, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 30, 551, 1092, 1456, 1663, 1623, 1676, 1587, 1798, 1898, 1799, 1453, 1957, 644, 2210, 281, 7254, 16774, 15160, 17118, 19362, 21795, 22140, 21917, 23356, 24622, 23248, 22432, 23053, 20738, 24381, 10669, 0, 1983, 110, 1082, 639, 960, 827, 847, 901, 786, 1003, 566, 2021, 3544, 2950, 3484, 3801, 4065, 4148, 4260, 4227, 4182, 4219, 4130, 3927, 3861, 4049, 3818, 3635, 3543, 3330, 2873, 2184, 1656, 523, 0, 55, 0, 15, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 276, 0, 984, 0, 9449, 20790, 21221, 23631, 23583, 25941, 25032, 25743, 25783, 26446, 26853, 27422, 27371, 26713, 27220, 26444, 27800, 25349, 30207, 14310, 0, 3117, 688, 3432, 3786, 4028, 4341, 4403, 4496, 4355, 4151, 4178, 4107, 4127, 4211, 4169, 4263, 4387, 4188, 4417, 4298, 4450, 4557, 4314, 4482, 4498, 4532, 4234, 4150, 4002, 4104, 3705, 3688, 1507, 0, 182, 0, 51, 0, 10, 0, 39, 0, 195, 0, 689, 0, 5565, 13113, 11388, 12682, 12055, 14342, 5546, 0, 653, 0, 193, 0, 54, 0, 170, 708, 1011, 1091, 1075, 1203, 1281, 1410, 1079, 748, 312, 0, 39, 0, 10, 0, 1, 0, 0, 0, 12, 0, 62, 0, 219, 0, 1793, 4282, 4181, 4679, 4501, 4836, 4906, 4797, 4794, 4585, 4060, 4436, 3718, 2846, 3159, 2734, 3377, 4525, 4663, 4997, 4950, 4613, 4682, 4317, 2410, 1258, 1442, 1348, 1429, 1537, 1480, 1593, 1682, 1813, 1768, 2458, 4236, 4767, 4660, 4700, 4689, 4676, 4727, 4500, 4064, 4164, 4071, 3771, 3344, 2968, 1763, 235, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 887, 0, 3151, 0, 20641, 20627, 0, 3857, 0, 1822, 533, 1124, 253, 0, 6, 32, 0, 245, 0, 884, 0, 7520, 19357, 20143, 22759, 24573, 26205, 26960, 26828, 27012, 23850, 25824, 11483, 0, 2509, 575, 1731, 1088, 1475, 1381, 1997, 2724, 3258, 3551, 3733, 4461, 4767, 4837, 4876, 5043, 5114, 5163, 5199, 5152, 5240, 5287, 5497, 5608, 5570, 5602, 5560, 5636, 5358, 4787, 4646, 4606, 4628, 4438, 4300, 3912, 3562, 1260, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 194, 0, 910, 0, 7333, 23432, 30566, 29528, 36790, 16379, 0, 2887, 314, 2322, 1942, 2069, 1527, 1895, 1077, 1916, 340, 2954, 0, 16469, 36143, 29004, 33121, 29262, 30892, 13262, 0, 3764, 2046, 3193, 2549, 2995, 3007, 3056, 3059, 3053, 3062, 3045, 3080, 2953, 2727, 2643, 2935, 3263, 3515, 3853, 4038, 4192, 4104, 4018, 4104, 4195, 3986, 3609, 1193, 0, 128, 0, 37, 0, 0, 47, 0, 252, 0, 875, 0, 7329, 17960, 15543, 16260, 15845, 15557, 15066, 15214, 15368, 14658, 13946, 14314, 13849, 14609, 13266, 15907, 7366, 0, 2657, 1697, 2230, 1674, 1894, 1771, 2020, 2169, 919, 304, 687, 112, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 4, 0, 137, 880, 1452, 1891, 2471, 2694, 2803, 2933, 3151, 3227, 3192, 3202, 3205, 3188, 3226, 3147, 3385, 3547, 3791, 4009, 3985, 4399, 4453, 3806, 3213, 3444, 3379, 3379, 2237, 975, 892, 1090, 1345, 2080, 3193, 3645, 4219, 4647, 4602, 4556, 4821, 4842, 4778, 4832, 4915, 4977, 4872, 4726, 4708, 4767, 4695, 4500, 4626, 4113, 3682, 3819, 3733, 3813, 3708, 3894, 3292, 2529, 2209, 1746, 606, 0, 67, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 92, 220, 163, 224, 131, 291, 0, 1010, 2165, 2044, 2029, 1710, 1740, 1977, 2078, 2117, 2026, 1882, 2068, 2401, 2544, 2596, 2576, 2599, 2541, 2431, 2662, 2388, 2322, 1976, 1620, 1690, 548, 0, 87, 0, 339, 1126, 1710, 2197, 2538, 2856, 3037, 3215, 3267, 3216, 3271, 3176, 3347, 3034, 3657, 1617, 0, 200, 0, 57, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 100, 0, 943, 2434, 2806, 3212, 3539, 2237, 857, 0, 1387, 0, 9904, 25243, 26922, 29474, 28436, 29034, 28601, 29074, 28318, 30618, 32815, 31923, 32079, 30119, 28452, 10519, 0, 2347, 581, 2176, 3275, 4210, 4440, 4368, 4328, 4374, 4241, 4064, 4087, 4226, 4334, 4421, 4479, 4502, 4366, 3977, 4012, 4185, 4151, 4153, 4165, 4164, 4036, 3890, 3804, 3724, 3657, 3632, 3678, 3580, 3769, 3419, 4119, 1822, 0, 226, 0, 64, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 13, 0, 44, 0, 465, 1638, 1914, 1984, 2163, 2288, 2618, 2560, 2696, 3017, 2815, 2858, 3051, 3084, 2901, 2907, 2822, 2751, 2778, 2715, 2941, 3138, 3166, 3163, 3166, 3161, 3172, 3145, 3254, 3367, 2820, 1793, 1342, 476, 0, 54, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 5, 1, 348, 1292, 584, 880, 0, 14875, 26450, 28530, 29079, 35789, 16866, 0, 3612, 541, 2147, 1040, 2028, 981, 1755, 0, 2375, 0, 16422, 36997, 30212, 33790, 27587, 30916, 13334, 0, 2196, 0, 1112, 295, 868, 243, 1921, 3709, 3310, 3494, 3393, 3664, 3595, 3606, 3785, 3733, 3655, 3610, 3519, 3375, 3378, 3335, 3092, 2921, 2241, 1865, 713, 0, 84, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 320, 0, 1113, 0, 8993, 20381, 16893, 18804, 15448, 4733, 0, 474, 0, 130, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 307, 0, 1061, 0, 9357, 25538, 25071, 28260, 29472, 30450, 31537, 31538, 31427, 31296, 31309, 31326, 31316, 31317, 30782, 27769, 28017, 11117, 0, 2517, 613, 2176, 2609, 3051, 3338, 2988, 2789, 2857, 2570, 2643, 2817, 2884, 2997, 3076, 3228, 3276, 3363, 3520, 3665, 3598, 3506, 3413, 3277, 2570, 1996, 2054, 653, 0, 66, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 0, 528, 0, 1857, 0, 14949, 34024, 29594, 32311, 30364, 30439, 28447, 28238, 27533, 28158, 27521, 25961, 8989, 0, 947, 0, 273, 0, 56, 0, 0, 0, 3, 0, 12, 0, 100, 91, 0, 13, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 382, 0, 1348, 0, 10818, 25212, 22403, 25700, 23018, 24812, 9333, 0, 1094, 0, 315, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 594, 1147, 1324, 1383, 1752, 1969, 1662, 1643, 1515, 1376, 1736, 1728, 1578, 1807, 1896, 1977, 1888, 1740, 1821, 2125, 2073, 2199, 1577, 1247, 646, 0, 88, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 170, 0, 884, 0, 3139, 0, 20588, 20803, 0, 4283, 0, 899, 0, 156, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 0, 381, 0, 1335, 0, 11405, 29672, 29548, 31572, 30832, 32072, 31696, 31622, 31520, 31059, 30098, 28744, 27053, 25534, 9092, 0, 1671, 318, 1245, 1003, 2198, 3164, 3449, 3575, 3783, 3898, 3722, 3728, 3747, 3678, 3589, 3544, 3596, 3497, 3683, 3340, 4024, 1780, 0, 221, 0, 63, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 189, 0, 668, 0, 7176, 19797, 24363, 28340, 28320, 29325, 29095, 29193, 29219, 29074, 28868, 29107, 24437, 26692, 11632, 0, 1373, 0, 391, 0, 92, 0, 1, 0, 7, 0, 173, 996, 1382, 1268, 1354, 1250, 1410, 1113, 2061, 2974, 2697, 2961, 2809, 2846, 2778, 2664, 2663, 2625, 2367, 1471, 317, 0, 24, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 137, 892, 1267, 1409, 576, 0, 70, 0, 21, 0, 15, 31, 97, 76, 174, 289, 252, 272, 259, 271, 253, 310, 378, 342, 219, 221, 31, 481, 1351, 1760, 1787, 1525, 1551, 1608, 1928, 2037, 1828, 615, 0, 67, 0, 19, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28246, 28894, 29871, 29592, 29574, 29422, 29624, 27441, 27776, 20452, 13905, 15694, 15118, 14862, 16180, 10997, 5185, 6593, 6244, 5719, 4473, 4768, 4249, 3637, 1201, 0, 131, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 27, 0, 76, 0, 1045, 4082, 1791, 0, 210, 0, 64, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 27, 0, 236, 563, 167, 36, 0, 249, 0, 2575, 2065, 8893, 14152, 10732, 14941, 19266, 35918, 15401, 0, 0, 15068, 35811, 26264, 28102, 27291, 28438, 27744, 27343, 27792, 28040, 27600, 27876, 28106, 28191, 28051, 27923, 27661, 27250, 27296, 27494, 27518, 27515, 27523, 27503, 27545, 27462, 27692, 27720, 27756, 27829, 27679, 28034, 27380, 26856, 26947, 27029, 26350, 25574, 25801, 25524, 25074, 25217, 25264, 25477, 25112, 25887, 26912, 26924, 26964, 27742, 24910, 21806, 17309, 4172, 0, 141, 172, 0, 3568, 10602, 7899, 5391, 4665, 4521, 4922, 4815, 4774, 4976, 4532, 5453, 2414, 0, 299, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 175, 0, 603, 0, 5070, 12533, 10668, 11707, 10221, 8437, 8115, 6743, 4447, 3923, 3635, 3306, 3698, 3089, 4229, 1892, 0, 235, 0, 18, 124, 0, 828, 0, 3096, 0, 20038, 18344, 0, 0, 15591, 34302, 15989, 5663, 0, 2112, 0, 7361, 13744, 11780, 13012, 11897, 13315, 10895, 18454, 25809, 22714, 23684, 23777, 23952, 24757, 26195, 28344, 31317, 31123, 33057, 30236, 35857, 16787, 0, 4841, 0, 17460, 35506, 29324, 31337, 28965, 25574, 21656, 22461, 21893, 21412, 21213, 21221, 20966, 20315, 20761, 20786, 21510, 23620, 24270, 24441, 24252, 24349, 24250, 24424, 24089, 24764, 22997, 23134, 19941, 18097, 9821, 0, 500, 0, 144, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 77, 0, 274, 0, 1797, 1797, 0, 272, 0, 59, 0, 0, 139, 0, 893, 1814, 9215, 14822, 15087, 14131, 20620, 26071, 34214, 16688, 0, 5196, 2413, 4078, 3184, 3632, 3560, 3889, 3453, 4090, 2083, 5105, 0, 15741, 34314, 28587, 31467, 29899, 30801, 30170, 30886, 29484, 31361, 29775, 36313, 16115, 0, 2925, 0, 3298, 0, 16933, 36975, 28690, 31133, 27863, 36511, 15848, 0, 2600, 3078, 0, 16450, 36058, 27969, 30646, 25419, 20450, 17715, 16860, 16548, 15798, 15196, 15038, 14298, 12844, 12443, 12022, 11735, 11946, 11602, 12217, 11101, 13319, 6038, 0, 694, 0, 199, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 215, 0, 814, 0, 6711, 15926, 20215, 24401, 33673, 15273, 0, 5040, 2720, 4848, 4207, 4772, 4673, 4918, 4930, 4920, 4592, 5241, 3730, 5877, 397, 16740, 33251, 28153, 30801, 29572, 30213, 29961, 29958, 30186, 29286, 28206, 28281, 28102, 28048, 28005, 27869, 27679, 27852, 27967, 28085, 28408, 28714, 28502, 28486, 28804, 29026, 29185, 29508, 29038, 28078, 28131, 28096, 28039, 28266, 28465, 28941, 28449, 28195, 25860, 24513, 25143, 23726, 21721, 19309, 17543, 16966, 17103, 16899, 17191, 16643, 17678, 15754, 19571, 7755, 477, 6841, 7106, 6250, 2329, 3998, 4704, 4508, 5191, 3305, 1420, 1323, 0, 215, 0, 54, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 594, 0, 2120, 0, 13833, 13681, 0, 4649, 1905, 4205, 3449, 4043, 3978, 4044, 3972, 3913, 4015, 3716, 3680, 1486, 4150, 0, 14486, 31819, 25768, 28316, 26900, 27610, 27338, 27321, 27595, 26588, 25716, 25761, 25067, 25451, 26122, 26641, 26861, 27089, 27423, 27414, 27437, 27596, 27648, 28257, 28333, 28463, 28403, 29344, 29690, 29107, 28810, 29037, 28849, 28226, 28367, 28652, 28070, 29660, 30388, 26944, 26018, 26410, 24836, 21708, 16641, 12826, 8740, 6170, 6965, 6483, 6908, 6374, 7290, 4583, 2585, 2477, 2089, 3312, 3431, 2872, 507, 0, 26, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 37, 0, 128, 0, 1528, 5901, 7786, 7316, 8174, 6533, 13726, 25104, 26446, 25638, 26406, 27600, 29877, 28008, 35579, 16060, 0, 2657, 377, 912, 2278, 0, 15009, 33388, 27637, 30232, 28364, 29350, 28856, 28880, 28854, 28843, 28844, 28854, 28828, 28884, 28705, 28593, 28764, 28798, 28885, 28889, 28806, 28806, 28717, 28783, 28674, 28804, 28933, 28694, 28702, 28312, 27998, 27960, 27563, 27259, 27790, 26905, 27280, 25377, 25822, 10013, 0, 1176, 0, 336, 0, 82, 0, 66, 0, 232, 0, 1863, 4253, 3454, 3985, 3463, 4182, 2904, 6755, 9203, 7581, 8596, 8042, 2946, 0, 332, 0, 91, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 242, 0, 858, 0, 7428, 18935, 18860, 18928, 25402, 28492, 35530, 16766, 0, 3957, 2268, 2396, 4676, 0, 16819, 36721, 30534, 33797, 31748, 33419, 30374, 28115, 28892, 28349, 28433, 28356, 28539, 28460, 28554, 28498, 28676, 28720, 28789, 28770, 28919, 29035, 28959, 29080, 29082, 28882, 29052, 28859, 29239, 28740, 29585, 23774, 11079, 8811, 3615, 0, 443, 0, 127, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 38, 0, 596, 2862, 3569, 4378, 5144, 5204, 5547, 5845, 2859, 487, 510, 0, 184, 0, 446, 0, 1427, 0, 12578, 33110, 25484, 29240, 32131, 27171, 25208, 25750, 25971, 29455, 14299, 0, 14681, 28909, 25106, 27016, 25878, 26639, 25980, 27306, 28443, 27859, 27958, 27646, 27392, 26931, 26545, 26361, 26081, 26097, 25936, 25902, 25994, 25604, 25973, 27028, 28262, 28588, 28486, 28727, 28534, 28639, 28395, 28449, 28849, 28796, 29450, 29431, 30470, 31587, 31037, 29557, 28653, 29092, 28110, 27939, 28226, 27968, 28275, 27761, 28671, 27025, 30350, 18575, 883, 360, 0, 126, 0, 8, 0, 0, 0, 1, 0, 9, 0, 35, 0, 255, 438, 301, 405, 357, 651, 287, 0, 35, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 35, 0, 310, 664, 4701, 15695, 25697, 25097, 33753, 16064, 0, 5800, 3238, 4916, 4151, 4604, 4502, 4558, 4627, 4754, 4810, 4487, 4101, 4064, 3824, 3674, 3724, 3683, 3734, 3656, 3758, 3417, 2552, 3360, 1744, 3990, 0, 14621, 33679, 28495, 29029, 28226, 28397, 28187, 28183, 28058, 27964, 28360, 27461, 29968, 25904, 35197, 16137, 0, 0, 13592, 33184, 26652, 29648, 27899, 27628, 28767, 26800, 31598, 13596, 0, 1668, 0, 466, 0, 28, 92, 0, 489, 0, 3828, 8447, 8232, 6621, 2565, 1078, 0, 363, 154, 0, 16, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 334, 0, 3043, 9046, 10904, 11362, 11369, 11075, 10522, 11023, 11238, 12980, 14080, 14337, 14221, 11361, 10370, 5262, 1273, 1187, 0, 202, 0, 48, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 40, 0, 135, 0, 1452, 5426, 6281, 6820, 6495, 6989, 3874, 1616, 1966, 4374, 3583, 11795, 21859, 22676, 26326, 26248, 27645, 28550, 29040, 29282, 29825, 30524, 30934, 31210, 30944, 31399, 30583, 32173, 27234, 23740, 26296, 25422, 25836, 17379, 15588, 16929, 18046, 18335, 22502, 10920, 0, 1253, 0, 356, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 124, 0, 433, 0, 3355, 6787, 4482, 4978, 3994, 3017, 3011, 3108, 3524, 2556, 4445, 627, 12802, 22599, 17737, 13988, 9708, 8479, 3644, 2876, 2089, 1021, 0, 126, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 157, 0, 547, 0, 4559, 11109, 9241, 10012, 10816, 14745, 14750, 17001, 21839, 23405, 25547, 26805, 23183, 20108, 17384, 9655, 7137, 8336, 8999, 9404, 9305, 9160, 8756, 8874, 7914, 5492, 4540, 3845, 2799, 4100, 1954, 0, 246, 0, 71, 0, 14, 0, 0, 0, 0, 0, 4, 0, 20, 0, 69, 0, 623, 1714, 1487, 1635, 2017, 2053, 2062, 1766, 2356, 1318, 0, 818, 3589, 7071, 9258, 11015, 11563, 12002, 12462, 13058, 14415, 15391, 16222, 16701, 16209, 17277, 12771, 7798, 7152, 5203, 5464, 5338, 6735, 6192, 4857, 5358, 5001, 5377, 4844, 5818, 2633, 0, 1844, 2829, 2763, 2966, 3145, 3042, 3298, 2609, 2004, 1375, 0, 3520, 14640, 21091, 17331, 7914, 4444, 1938, 135, 2201, 1832, 2756, 1190, 0, 65, 0, 6, 17, 0, 105, 0, 1021, 3239, 4086, 4380, 4840, 5293, 5170, 5198, 5243, 5106, 5413, 4357, 2749, 939, 0, 88, 0, 0, 230, 345, 789, 1855, 1922, 2100, 2101, 2924, 4213, 2555, 314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 232, 1813, 4228, 5072, 4808, 5066, 4696, 5312, 4138, 7957, 11701, 9716, 11454, 6017, 71, 184, 0, 66, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 52, 0, 188, 0, 1379, 2408, 1709, 1934, 2396, 3512, 3274, 2915, 3974, 4171, 4117, 2102, 0, 117, 0, 0, 440, 723, 2268, 4388, 4639, 4634, 3984, 1313, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 114, 0, 400, 0, 3278, 7799, 6982, 7941, 7847, 8725, 7721, 10850, 13581, 10742, 16475, 19671, 18221, 18858, 17800, 17377, 17592, 17616, 18744, 13171, 3615, 5519, 10141, 10675, 10292, 9694, 10115, 10573, 10441, 10512, 10464, 10503, 10507, 9661, 3423, 0, 949, 155, 28, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 51, 0, 235, 0, 1251, 467, 5487, 11977, 16407, 23321, 24567, 25379, 26023, 27241, 29481, 30340, 31314, 32582, 32075, 31723, 31235, 31451, 31249, 31528, 31060, 31973, 28890, 24602, 22450, 18579, 18230, 18450, 17682, 16721, 16504, 15009, 14405, 12995, 11334, 12249, 8707, 2686, 67, 29, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 36, 50, 1199, 1141, 2317, 3277, 3659, 4744, 4411, 4487, 4618, 4235, 5077, 2251, 0, 279, 0, 79, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 53, 0, 176, 0, 1489, 3578, 2147, 3157, 2676, 1540, 2159, 2861, 1143, 0, 0, 549, 0, 5292, 13149, 12478, 13024, 14064, 13246, 15033, 6674, 0, 828, 0, 220, 0, 0, 138, 144, 1014, 1773, 1530, 1445, 1017, 1077, 1261, 1301, 1311, 1277, 1344, 1219, 1469, 650, 0, 80, 0, 22, 0, 14, 0, 48, 0, 136, 0, 1730, 4515, 3202, 4617, 689, 5239, 15984, 14961, 16243, 21597, 25367, 26862, 27130, 26911, 26499, 25801, 23903, 20123, 18598, 18133, 18235, 19001, 19287, 17590, 16869, 15407, 13840, 14491, 13870, 14735, 13297, 16070, 7088, 0, 834, 0, 1440, 401, 0, 40, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 491, 663, 951, 2261, 2706, 4210, 5857, 6332, 5859, 5336, 5830, 5412, 5585, 5560, 5027, 4929, 4897, 4989, 4807, 5150, 4473, 6462, 6623, 3978, 3837, 4151, 3244, 3099, 3698, 4332, 4719, 1999, 284, 0, 10, 0, 0, 10, 0, 75, 99, 0, 100, 0, 314, 0, 2139, 2092, 0, 306, 0, 49, 28, 0, 582, 1310, 702, 1436, 2141, 2077, 2139, 2087, 2144, 2062, 2212, 1695, 923, 776, 208, 0, 18, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 18, 0, 62, 0, 697, 2686, 3483, 3738, 3773, 3916, 3724, 4063, 1641, 0, 192, 0, 55, 0, 11, 0, 0, 0, 0, 3, 0, 39, 0, 362, 1002, 2248, 1020, 5882, 9770, 7157, 5982, 4484, 4804, 4214, 3444, 3156, 2777, 2903, 3333, 2965, 2391, 1759, 1146, 266, 0, 22, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 34, 0, 134, 0, 1035, 2491, 4233, 3395, 2010, 4149, 7376, 11064, 14194, 15596, 16779, 18514, 18459, 18116, 20589, 20147, 19912, 19419, 19425, 21476, 21463, 21927, 19397, 18794, 17565, 16035, 14851, 14029, 14009, 13892, 13633, 14294, 12991, 15639, 6922, 0, 859, 0, 246, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 66, 0, 306, 0, 1393, 0, 8807, 17664, 15583, 18046, 17929, 18944, 19735, 19145, 21651, 24039, 23365, 23626, 23620, 23345, 24504, 25474, 24808, 25484, 23978, 21478, 19954, 21518, 19768, 20072, 24272, 21980, 25421, 14635, 3013, 6724, 2320, 0, 4300, 2645, 0, 335, 0, 103, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 200, 0, 699, 0, 5784, 13786, 11895, 12375, 12035, 11809, 13333, 16274, 17591, 18410, 19097, 19828, 19180, 20742, 21556, 22010, 23512, 24802, 26468, 26578, 27274, 27319, 28312, 29597, 30434, 29912, 28814, 29426, 30870, 31911, 30947, 31923, 29374, 31156, 15825, 505, 0, 10251, 21294, 17713, 19801, 18092, 20107, 16936, 24077, 12977, 0, 1409, 0, 891, 3157, 2830, 7670, 11990, 5299, 2790, 3402, 3788, 6532, 5969, 12185, 19997, 22061, 23564, 20789, 13864, 10339, 11727, 11149, 11029, 10229, 10019, 5024, 2878, 3033, 647, 262, 0, 39, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 71, 0, 222, 0, 3075, 5438, 3651, 5225, 1233, 5469, 14403, 12904, 19277, 26289, 27818, 27676, 29292, 24888, 18275, 18702, 18030, 18515, 17978, 18779, 17398, 20112, 11300, 2963, 5837, 4248, 4567, 4151, 1645, 0, 183, 0, 52, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 62, 0, 235, 0, 1644, 2835, 3581, 2939, 879, 1306, 1617, 500, 2833, 0, 13962, 30476, 24480, 26823, 18833, 16324, 12337, 6939, 7873, 7286, 3158, 0, 320, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 304, 0, 1063, 0, 8491, 18564, 14432, 18957, 21814, 20053, 15305, 15139, 15610, 18483, 19317, 25280, 31834, 30884, 32395, 30464, 27880, 24504, 13318, 7993, 9081, 8272, 8144, 7817, 7180, 4849, 1870, 0, 61, 0, 17, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 47, 0, 193, 0, 1390, 3077, 7626, 13357, 15781, 17070, 17057, 16266, 15762, 16624, 15430, 13131, 13547, 15334, 14542, 15407, 8053, 2322, 4180, 3885, 4604, 4956, 5243, 5330, 5221, 5385, 5881, 5857, 5744, 5487, 4802, 3653, 1035, 0, 101, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 20, 0, 97, 0, 322, 0, 2888, 7922, 6826, 9563, 10197, 9007, 10012, 9728, 10888, 11126, 11108, 9760, 9438, 7117, 6605, 4905, 10697, 16934, 16955, 20941, 22128, 24583, 27293, 29918, 30316, 30763, 30894, 30987, 30716, 31269, 30215, 32357, 25090, 15415, 12293, 9336, 9772, 8502, 8153, 7323, 5495, 4174, 3493, 3246, 2885, 2773, 1254, 0, 158, 0, 43, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 158, 477, 1835, 962, 5167, 10071, 9790, 10475, 10133, 10348, 10180, 10365, 10025, 11620, 15569, 12009, 7850, 8291, 8947, 9660, 10035, 10370, 10594, 10116, 9106, 8011, 6747, 6896, 6583, 6086, 5749, 4872, 5738, 2423, 0, 294, 0, 84, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 0, 370, 0, 1304, 0, 10915, 27192, 26155, 27785, 27515, 28944, 26540, 25427, 23119, 22610, 22659, 22991, 22004, 21243, 21987, 20817, 20475, 19753, 19761, 19555, 19298, 19225, 18757, 17821, 17634, 17476, 16628, 12636, 10868, 12694, 11325, 9619, 3188, 0, 349, 0, 101, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 130, 0, 450, 0, 3432, 6626, 4199, 6090, 5053, 1463, 0, 1085, 3127, 4107, 6660, 9248, 10110, 10665, 12122, 12112, 11790, 13148, 14061, 13581, 10033, 2729, 0, 259, 0, 73, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 104, 0, 346, 0, 3144, 8727, 6790, 8414, 9434, 8985, 6673, 5944, 3693, 6328, 13606, 17574, 20540, 21582, 19817, 16586, 11670, 7902, 8840, 8706, 8182, 9681, 4326, 0, 535, 0, 153, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 0, 92, 295, 322, 261, 577, 2804, 3816, 3801, 3398, 4336, 2331, 9263, 17683, 16775, 17817, 18013, 17019, 17538, 13146, 9150, 8924, 9811, 4513, 0, 567, 0, 156, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 149, 0, 531, 0, 4247, 10052, 10194, 7232, 716, 18, 0, 2, 85, 229, 0, 1441, 0, 5000, 0, 22866, 21195, 0, 11166, 9357, 11385, 9915, 7570, 6251, 5062, 3811, 4060, 1161, 0, 106, 0, 34, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 0, 158, 659, 518, 802, 0, 4002, 10840, 12173, 13472, 14129, 15230, 15290, 15951, 16604, 17162, 16242, 13773, 13419, 7399, 1044, 519, 0, 97, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 13, 0, 27, 502, 4908, 5733, 6682, 11241, 8609, 1983, 0, 1012, 1835, 4558, 6486, 7988, 9383, 9858, 9896, 9755, 9875, 9794, 9893, 9733, 10015, 9454, 11339, 13539, 12872, 11888, 10826, 10515, 9829, 9399, 8741, 8069, 8280, 6749, 1748, 0, 153, 0, 44, 0, 10, 0, 0, 0, 0, 0, 0, 27, 0, 131, 0, 457, 0, 3718, 8442, 7106, 11287, 14954, 15435, 14596, 14421, 14348, 14575, 14107, 14989, 13209, 19237, 26504, 25589, 26607, 26873, 26905, 25026, 20788, 16907, 11798, 10093, 4166, 0, 510, 0, 141, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 54, 0, 179, 0, 1518, 3443, 853, 0, 107, 980, 1152, 1152, 1104, 3504, 5863, 12850, 17958, 18624, 20353, 21910, 21201, 18547, 17094, 16906, 9082, 1240, 1146, 0, 210, 0, 45, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 135, 0, 495, 0, 3968, 9704, 11533, 14497, 15527, 20109, 13547, 1840, 3892, 10457, 12599, 14259, 14268, 12075, 11592, 11620, 10962, 10941, 10853, 10624, 10818, 10498, 11071, 10032, 12093, 5349, 0, 664, 0, 190, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 0, 0, 998, 8574, 12382, 11983, 7243, 3557, 7770, 6567, 3095, 1068, 2105, 3101, 6367, 6434, 6657, 10555, 11470, 12138, 11916, 11994, 12007, 11909, 12136, 11346, 10353, 10435, 9936, 10101, 10110, 10256, 8925, 7043, 2406, 0, 269, 0, 75, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0);

--    type t_reg_datos is array (0 to 16391) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (20281, 19442, 16957, 15142, 15412, 15158, 15446, 15015, 15796, 13576, 13213, 14746, 14148, 13681, 14541, 16329, 16067, 17112, 17673, 17879, 17338, 16618, 17513, 17677, 18974, 19412, 19299, 20713, 20716, 21630, 19675, 17264, 17171, 15561, 14850, 14784, 14268, 13055, 12547, 12652, 15122, 16961, 15195, 15539, 15896, 16354, 18070, 17031, 15867, 16308, 15920, 16433, 15532, 18360, 21149, 20358, 20118, 20773, 18637, 15919, 16950, 15582, 14798, 14490, 13714, 12949, 12545, 12596, 14971, 15943, 14995, 15356, 15244, 15672, 15149, 16057, 12456, 12160, 14705, 14746, 17536, 19683, 20632, 19339, 18951, 18961, 18166, 16160, 14775, 13998, 13819, 14098, 13968, 14087, 13927, 14190, 13695, 15172, 15826, 15349, 15793, 15411, 15282, 15425, 13628, 10017, 13746, 17765, 18410, 19097, 18160, 18291, 18266, 18194, 16299, 14385, 14564, 14430, 14794, 15266, 14333, 13756, 13479, 13309, 14106, 14906, 15300, 15144, 15461, 16010, 15456, 16309, 13637, 10992, 11725, 11282, 11449, 11483, 11226, 11807, 10600, 14305, 16406, 15236, 13275, 13058, 15040, 13489, 14385, 13898, 13520, 14624, 14786, 15443, 16125, 15897, 16159, 16090, 16773, 16294, 17475, 13735, 13670, 18340, 18214, 19152, 18688, 18990, 19240, 18986, 18450, 16352, 15067, 14897, 14771, 13998, 13388, 13457, 13339, 13298, 13285, 13327, 13245, 13388, 13092, 14315, 16772, 14728, 11917, 10636, 15085, 21140, 22611, 22406, 19945, 18489, 18989, 17788, 16992, 14503, 12555, 13098, 12361, 12425, 12993, 13356, 13007, 12966, 16652, 20103, 14402, 12960, 15909, 16334, 17999, 14797, 12790, 12737, 15005, 21705, 24848, 24482, 20347, 18059, 18770, 18263, 18819, 18002, 19501, 14603, 9666, 13565, 13866, 12085, 13051, 17623, 19252, 14209, 14067, 15731, 15216, 18963, 15817, 11225, 14981, 17980, 20281, 24541, 22807, 20467, 19093, 17833, 17734, 17626, 14109, 11981, 12690, 12902, 14158, 12030, 12482, 11230, 12450, 15248, 18058, 13732, 10762, 13912, 12626, 13377, 12833, 13384, 12527, 15303, 19022, 17438, 14309, 12046, 12024, 11579, 10825, 10179, 9118, 8125, 2635, 0, 255, 65, 1114, 3226, 7181, 4937, 4904, 5229, 2274, 2739, 3468, 3943, 3801, 7301, 6678, 7174, 10900, 8869, 8498, 8904, 9335, 9643, 7035, 3477, 966, 593, 639, 616, 637, 614, 646, 432, 0, 920, 1607, 2215, 1551, 3975, 8143, 8214, 10267, 9741, 7938, 10131, 10187, 7457, 5714, 6561, 8137, 8270, 7601, 2265, 0, 225, 0, 67, 0, 14, 0, 26, 0, 137, 0, 490, 0, 3741, 7569, 6772, 8447, 7694, 8055, 7896, 7942, 7960, 7852, 8708, 10921, 4059, 0, 455, 0, 149, 0, 108, 0, 273, 0, 1795, 1923, 0, 581, 0, 2464, 5584, 6427, 7625, 6219, 6980, 7178, 7515, 9055, 9759, 8363, 8337, 3322, 0, 396, 0, 113, 0, 22, 0, 0, 5, 0, 25, 0, 85, 0, 1129, 5119, 7333, 7720, 7425, 6328, 7226, 7642, 8519, 10360, 9287, 10455, 4203, 0, 502, 0, 146, 0, 29, 0, 0, 0, 0, 22, 0, 107, 0, 365, 0, 3117, 7916, 6425, 6725, 6224, 6632, 7095, 7462, 9068, 9327, 9414, 9186, 9628, 8807, 10461, 4833, 0, 1652, 748, 0, 56, 0, 0, 79, 0, 1299, 5605, 7450, 7420, 8089, 7137, 7347, 7928, 7175, 8053, 8066, 7902, 6757, 1869, 0, 216, 0, 165, 0, 1621, 6307, 2332, 684, 2183, 0, 958, 48, 3849, 7098, 6110, 6637, 6305, 6562, 6266, 7096, 8173, 7923, 8830, 8909, 8653, 7891, 6772, 2250, 0, 0, 1635, 7379, 8126, 8533, 10605, 7486, 1583, 3259, 5942, 7265, 9388, 10075, 10243, 10946, 13124, 15126, 11046, 7483, 9598, 10056, 10725, 9051, 7840, 7345, 7244, 6372, 3654, 2900, 3028, 2991, 2975, 3060, 2833, 3762, 6458, 10692, 11310, 10331, 10642, 12155, 15508, 15761, 16054, 13437, 11339, 14072, 13996, 13475, 12873, 11615, 12032, 12772, 10522, 7813, 8735, 8864, 8034, 11356, 15652, 11520, 7766, 9196, 10968, 13339, 11543, 9800, 11402, 15953, 17335, 17562, 17249, 15480, 16118, 15775, 15985, 15834, 16004, 15238, 12837, 13847, 12237, 10779, 9816, 11283, 14596, 15024, 13224, 8358, 11357, 13157, 13102, 14028, 11838, 15129, 18273, 18704, 20247, 19379, 17872, 16548, 16950, 16816, 14881, 15317, 15546, 15735, 14612, 14881, 14038, 11290, 11287, 13466, 14409, 16901, 14288, 10132, 11380, 10918, 10863, 11461, 9962, 15185, 20963, 20440, 20258, 19894, 19252, 16721, 17812, 14863, 14061, 16449, 16516, 15066, 13806, 13506, 10511, 11441, 14931, 16351, 18347, 16891, 14023, 17214, 17828, 17517, 14797, 11401, 17224, 20947, 20630, 21565, 21323, 20805, 20329, 19229, 16600, 14057, 14093, 14225, 14196, 14227, 14176, 14268, 14082, 14738, 16248, 17976, 16379, 13947, 16160, 16820, 17745, 15421, 9689, 14072, 19190, 19611, 20900, 20795, 20884, 20767, 19269, 18155, 15030, 13536, 14480, 14349, 14608, 14567, 15113, 14789, 13605, 15000, 18023, 18708, 18917, 16311, 16784, 19585, 18798, 20182, 16139, 12803, 13937, 13105, 14026, 12562, 17046, 21469, 18214, 15494, 14608, 14335, 15595, 15708, 14321, 15321, 15338, 14314, 14613, 17024, 18941, 18795, 16204, 16422, 19190, 18850, 20022, 15168, 11334, 17152, 19513, 19939, 21029, 20792, 20773, 20717, 17569, 16641, 16440, 16247, 16519, 16473, 15031, 14039, 14823, 14592, 14811, 14553, 14947, 14206, 16551, 18821, 19041, 18723, 14112, 11088, 15502, 19163, 18715, 19994, 20587, 20987, 19883, 17590, 16950, 15847, 14356, 15459, 16560, 15901, 15070, 13276, 11730, 13861, 15860, 17149, 18856, 18175, 17988, 18517, 18748, 19746, 14428, 10815, 16516, 19356, 19377, 19850, 19812, 19905, 19801, 19949, 19712, 20165, 18572, 16401, 17048, 14936, 15206, 15173, 14653, 16057, 17998, 18218, 15804, 16545, 18333, 18704, 19847, 15051, 9722, 16100, 19637, 19678, 20378, 19918, 20081, 19661, 18705, 16859, 15487, 14896, 14466, 14827, 15808, 15330, 17227, 14345, 13736, 17507, 17594, 18899, 18851, 18930, 18910, 18884, 18956, 18811, 19247, 19599, 20003, 20339, 20718, 20920, 20182, 19225, 17674, 17306, 17460, 17100, 16879, 16271, 16435, 16475, 16062, 16113, 17085, 18384, 20138, 21258, 20815, 20745, 19765, 21504, 18647, 15977, 18963, 20229, 21507, 22091, 22165, 21312, 20594, 20249, 20086, 18347, 17225, 17521, 17407, 17412, 17514, 17241, 18278, 19862, 20198, 21729, 23169, 23408, 22883, 21507, 22092, 22299, 21487, 20842, 20550, 21584, 21844, 21899, 21064, 20738, 20364, 18778, 17499, 17717, 17025, 16836, 16756, 16831, 17719, 16325, 15754, 16647, 16994, 18597, 19550, 18348, 18831, 18222, 20358, 15940, 11093, 12523, 11935, 12015, 12410, 11312, 15033, 17790, 16113, 16788, 13767, 13143, 15471, 15399, 15222, 14088, 12380, 10638, 13166, 15917, 16319, 17270, 16409, 16357, 15903, 18089, 13695, 11388, 11669, 13521, 17531, 18329, 17603, 16121, 17036, 15898, 16002, 13961, 12099, 13014, 14431, 14699, 15430, 13642, 11681, 12209, 12095, 11880, 12510, 11113, 15743, 20361, 20093, 19120, 17094, 20220, 20611, 19873, 20153, 20818, 20987, 20723, 20660, 18043, 16835, 16638, 17312, 18536, 18256, 18722, 18593, 18417, 18077, 19014, 20006, 20503, 21940, 21918, 21666, 21331, 21651, 21623, 20151, 20580, 20505, 19919, 19328, 19539, 20230, 19988, 20130, 20013, 20156, 19934, 20203, 17684, 16194, 16945, 17566, 16462, 16662, 18657, 19169, 20838, 20501, 20893, 20445, 20656, 20855, 19221, 19501, 19071, 18286, 17645, 18226, 19728, 19857, 20516, 19829, 17174, 15080, 15992, 16471, 15062, 14414, 13557, 13869, 14218, 15119, 17115, 18691, 18914, 18580, 18709, 18616, 18724, 18551, 18863, 18133, 18364, 15830, 13589, 15120, 14713, 15246, 16053, 15521, 15152, 15590, 15633, 15438, 15363, 14548, 13330, 13065, 14661, 15036, 17719, 18408, 18015, 20394, 20470, 21159, 20305, 19571, 19192, 19492, 19246, 16803, 17856, 18577, 18772, 18754, 18662, 19031, 18623, 19072, 18914, 18941, 19025, 18804, 19273, 17786, 16972, 18806, 19569, 20623, 20650, 19968, 19779, 18803, 18441, 17596, 18267, 19323, 17268, 17503, 18558, 18968, 20062, 19570, 19947, 19936, 20530, 20483, 18232, 17304, 16281, 16731, 17839, 19169, 17754, 18701, 19890, 21362, 20445, 19595, 20930, 19705, 20613, 20545, 20641, 20571, 20645, 20532, 20743, 20109, 20049, 21585, 21041, 21547, 20597, 19792, 19844, 18925, 18633, 19976, 20369, 18756, 19835, 20773, 22396, 21882, 21399, 22636, 21728, 21979, 22119, 21897, 22238, 21543, 20891, 20668, 20976, 21683, 21640, 21151, 22192, 21458, 19742, 20137, 19120, 18131, 18930, 19300, 19174, 19329, 19066, 19537, 18628, 21372, 22940, 22010, 23210, 22055, 23772, 24015, 22753, 22965, 22504, 22424, 22446, 22208, 22751, 22751, 22768, 21805, 21795, 21022, 19172, 20004, 20124, 21045, 22316, 21595, 20749, 20764, 22691, 23159, 21718, 21988, 23110, 22205, 23220, 24502, 23425, 24121, 23879, 23631, 23717, 23640, 23736, 23589, 23865, 22931, 21683, 21929, 22501, 21997, 21229, 22531, 23140, 22670, 22846, 22199, 22367, 21840, 21632, 22843, 23079, 22151, 22119, 23459, 23930, 24182, 22964, 22752, 22965, 22415, 23357, 23692, 22440, 22035, 21641, 21550, 22266, 22083, 22797, 23654, 23153, 22047, 22150, 22662, 22496, 22577, 22540, 22546, 22567, 22583, 23494, 24453, 24971, 23851, 23081, 23220, 22914, 22993, 22507, 22303, 22661, 22018, 21586, 22611, 21584, 23130, 24542, 22856, 22155, 22283, 22374, 23379, 22852, 22123, 23380, 22802, 23146, 23936, 24669, 25235, 24608, 24078, 23536, 22986, 22137, 21445, 22548, 23201, 23025, 23122, 23049, 23124, 23024, 23173, 22101, 20162, 20176, 21106, 21454, 21176, 21326, 21634, 21672, 22184, 22296, 23203, 23916, 23891, 22567, 21314, 20336, 20060, 20993, 21167, 21249, 21164, 21288, 20632, 20546, 20042, 21467, 23147, 21406, 19880, 19827, 20252, 21058, 20462, 19998, 21131, 20520, 19988, 20137, 20057, 20108, 20072, 20112, 19919, 19052, 18484, 18284, 18523, 18777, 17661, 17295, 16575, 17365, 18433, 20520, 20103, 17864, 18706, 19168, 20000, 20184, 19944, 19534, 18360, 19710, 21108, 21214, 22027, 21600, 21043, 19431, 18358, 17862, 17880, 17746, 17216, 17310, 16892, 16206, 16297, 16576, 16563, 16549, 16614, 16468, 16755, 16172, 17987, 19090, 18354, 18165, 19711, 19827, 18805, 20217, 19896, 18950, 18080, 17749, 17409, 17081, 16151, 15824, 14641, 14602, 15526, 15361, 14517, 15111, 14635, 16489, 17884, 16678, 17309, 17983, 19085, 18465, 18285, 17317, 18171, 18945, 18097, 19197, 19909, 19158, 18823, 18776, 19008, 18520, 19528, 16160, 12615, 13650, 13447, 14573, 14711, 14870, 16331, 16913, 16365, 16170, 17020, 18034, 17324, 16363, 15948, 17105, 18052, 18041, 18207, 18521, 17600, 16925, 16203, 15367, 15007, 14359, 14672, 14163, 13598, 13649, 13702, 14018, 14805, 14622, 14979, 15816, 15701, 16476, 17066, 16907, 16963, 16981, 16876, 17154, 17083, 18845, 19087, 17665, 18386, 16635, 15991, 14861, 14353, 15129, 14246, 14322, 13996, 14161, 14402, 14842, 14656, 14770, 15819, 15910, 16360, 15903, 16336, 15398, 11657, 14541, 18052, 17135, 17478, 17790, 18248, 17843, 17523, 16147, 15325, 13228, 11507, 13367, 13622, 13703, 13553, 13815, 13306, 14774, 14717, 12966, 13157, 14140, 15909, 16019, 16663, 13971, 15076, 18813, 18232, 19076, 18629, 17955, 17800, 17424, 17025, 15942, 15830, 15862, 15995, 15034, 14499, 14539, 14189, 14973, 15755, 14871, 12697, 12235, 12300, 13476, 15618, 15720, 16529, 14521, 15926, 18815, 17862, 18357, 18067, 18263, 18083, 18275, 17001, 15817, 14654, 13660, 14348, 13337, 14686, 12378, 12461, 15777, 15419, 13850, 13204, 14400, 14703, 16901, 17308, 14988, 12878, 16271, 18966, 18395, 19010, 18285, 17857, 17803, 17834, 18601, 17024, 15687, 16041, 16588, 16871, 15002, 14425, 14693, 15134, 15743, 15512, 15672, 15517, 15720, 15354, 16740, 18778, 15919, 16679, 19339, 18116, 17912, 18139, 17935, 17791, 17812, 18008, 16714, 15010, 16251, 16784, 16585, 15701, 15116, 14448, 15071, 16740, 17171, 17107, 16663, 17124, 17614, 18261, 18404, 18764, 18443, 18376, 19021, 17875, 17218, 17698, 17424, 17199, 17121, 17164, 17100, 17214, 17007, 17419, 16079, 14938, 16210, 16952, 17556, 16829, 15975, 16347, 17029, 17410, 17629, 18323, 18434, 18004, 18807, 18448, 17900, 18317, 18301, 18236, 17581, 18060, 17616, 16960, 17066, 17034, 16113, 15246, 15743, 16570, 15383, 15784, 17132, 16029, 16049, 16903, 17405, 17475, 17765, 17661, 17717, 17680, 17716, 17660, 17860, 18320, 18572, 18097, 18032, 17589, 15921, 14980, 15054, 15033, 15140, 16526, 13353, 10618, 15439, 16819, 16681, 16398, 15656, 16736, 16983, 17792, 19086, 17095, 16842, 18838, 17748, 17796, 17886, 18139, 18496, 18178, 18269, 17407, 16940, 17342, 17239, 15912, 14954, 15222, 15109, 15136, 15184, 15029, 15598, 16415, 17089, 17636, 18048, 18791, 17820, 17721, 18177, 17058, 16788, 17769, 18406, 18055, 17898, 16939, 16416, 15497, 13603, 14502, 14278, 15185, 14619, 13733, 15205, 15537, 16479, 15931, 15313, 16704, 17438, 17835, 17097, 15877, 14594, 16431, 18264, 17037, 17322, 17181, 17167, 17351, 16930, 17808, 15045, 12894, 12793, 13546, 14110, 12176, 10790, 13836, 17425, 15847, 15136, 13414, 13862, 14867, 15067, 16260, 16048, 14548, 16361, 18112, 17303, 17213, 17507, 17628, 17411, 17414, 16276, 16212, 15062, 13954, 12458, 12290, 12812, 10822, 13126, 16335, 17302, 15525, 14296, 14607, 14526, 14441, 14723, 14086, 16224, 18269, 17334, 17375, 17076, 17724, 17604, 17275, 17266, 17348, 15843, 13985, 15081, 14478, 14844, 13655, 13911, 16738, 16893, 17977, 16885, 15335, 16273, 16740, 17285, 18492, 18491, 18002, 18105, 18475, 18117, 17811, 17633, 17935, 17581, 17696, 16669, 16406, 17296, 16970, 17139, 17051, 17086, 17081, 17209, 18090, 16558, 14379, 13579, 15512, 17210, 17202, 14957, 15364, 18369, 18080, 18562, 18350, 18228, 18611, 18019, 17835, 17374, 16867, 16650, 15941, 16107, 16678, 16272, 16083, 15410, 16690, 17332, 16519, 15884, 15363, 15054, 16548, 17279, 16660, 15713, 16437, 18564, 17841, 18216, 17994, 18153, 17990, 18223, 17192, 16175, 16085, 16095, 16032, 16423, 16627, 16036, 15876, 16265, 16877, 16682, 16139, 16147, 16167, 17701, 18223, 17249, 18594, 19373, 19811, 19952, 19605, 19665, 18873, 18260, 17844, 18564, 17596, 16249, 16597, 16242, 16554, 16483, 15998, 15924, 15965, 15802, 15844, 15857, 15783, 15947, 15608, 16681, 17591, 17964, 19396, 19880, 19763, 19132, 19458, 19256, 17883, 17782, 18291, 17106, 15893, 17079, 17446, 17765, 17078, 16026, 15909, 16355, 17300, 17428, 16956, 17340, 18382, 18010, 18212, 18405, 18846, 19310, 19805, 19449, 19257, 18809, 18539, 18562, 17917, 17967, 17933, 17914, 17995, 17824, 18173, 17054, 15949, 15693, 15648, 16941, 17157, 16957, 17892, 18463, 18091, 18349, 18712, 18970, 18792, 18313, 18964, 19168, 19168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 75, 0, 327, 0, 2770, 6270, 5629, 0, 10661, 24447, 17811, 19006, 19355, 19646, 19980, 20235, 20679, 21353, 21611, 21753, 21756, 21986, 22034, 22426, 22159, 21898, 22147, 21543, 22148, 22492, 24410, 26015, 25737, 25488, 26324, 24583, 28178, 16344, 4833, 8428, 6593, 6552, 7611, 8549, 4108, 632, 3266, 2319, 0, 324, 0, 91, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 166, 0, 576, 0, 8443, 8730, 7098, 22821, 26982, 26424, 26509, 26703, 26127, 27444, 22951, 18922, 21343, 20781, 21230, 21519, 22905, 23671, 23448, 23399, 23198, 22542, 22695, 22738, 25128, 27074, 25322, 25960, 23176, 24912, 12790, 3700, 8316, 7956, 8945, 4867, 5206, 5986, 5111, 3746, 3574, 1577, 0, 196, 0, 54, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 174, 0, 554, 0, 5199, 12994, 1916, 5313, 22010, 27454, 27960, 27468, 27463, 26800, 23059, 21250, 21225, 20984, 19712, 19163, 19173, 18763, 18107, 17169, 17859, 18692, 20813, 21527, 24366, 26665, 25340, 28365, 30588, 30068, 30126, 30475, 29568, 31511, 25536, 21279, 16147, 7399, 4923, 311, 75, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 294, 0, 1040, 0, 8931, 21965, 16425, 12226, 21437, 30903, 29576, 30227, 29736, 28170, 26731, 27242, 26845, 27329, 26553, 28018, 23431, 19770, 21580, 21012, 21954, 21957, 22336, 22771, 24640, 27616, 28873, 26922, 28504, 28949, 29880, 23396, 14565, 7326, 2179, 3496, 1657, 1788, 1404, 1757, 811, 0, 236, 266, 120, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 35, 0, 93, 765, 9327, 12286, 13119, 24147, 29733, 30656, 31220, 30030, 32372, 27234, 37030, 10691, 13284, 36475, 33755, 17856, 0, 4576, 122, 1833, 1801, 1645, 1730, 3958, 2798, 2471, 2253, 5341, 0, 18031, 31694, 23601, 25727, 22468, 23920, 23467, 23181, 24253, 22038, 26537, 11743, 0, 1458, 0, 417, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 216, 0, 778, 0, 5941, 12045, 11512, 15774, 18464, 26572, 30758, 31092, 31141, 31175, 30307, 29069, 26263, 24898, 24061, 22585, 22786, 22689, 22605, 22975, 22125, 23882, 22341, 33055, 17070, 0, 4778, 1280, 4412, 1885, 5695, 0, 16400, 34338, 21858, 22097, 19843, 21733, 9119, 0, 1501, 0, 328, 0, 3008, 5137, 5295, 5962, 6283, 6140, 6914, 2769, 0, 322, 0, 59, 268, 2222, 3583, 3399, 3354, 3273, 3442, 3125, 3762, 1666, 0, 206, 0, 59, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 353, 0, 1275, 0, 9351, 17532, 18463, 30582, 30982, 31375, 27701, 24183, 20862, 19427, 20510, 19734, 19898, 20062, 21080, 21131, 22754, 25385, 26120, 26485, 26731, 28236, 27219, 29519, 28584, 36394, 15409, 201, 545, 17031, 32934, 26218, 30123, 23444, 23860, 21479, 18098, 6727, 657, 2318, 1469, 1997, 1594, 2053, 876, 0, 111, 0, 31, 0, 1, 5, 0, 41, 0, 144, 0, 1311, 4248, 4409, 4212, 2587, 8190, 4959, 0, 678, 0, 194, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 173, 0, 558, 0, 4903, 13632, 10760, 12193, 4752, 14757, 26826, 24124, 22492, 17886, 20167, 19542, 19687, 19751, 19643, 19596, 19744, 19678, 19460, 19679, 21084, 21918, 21980, 22161, 22032, 22210, 21909, 22467, 21345, 24946, 28216, 29992, 30717, 32290, 24487, 20713, 13511, 2448, 2781, 6145, 10501, 8753, 5454, 2112, 4543, 5401, 5458, 5418, 4968, 5741, 2480, 0, 305, 0, 83, 0, 0, 34, 0, 152, 0, 1194, 2653, 2411, 1643, 111, 23, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 336, 0, 1172, 0, 9465, 21532, 17930, 20160, 19409, 20137, 19972, 20464, 21598, 22190, 22062, 22117, 22121, 20881, 21115, 22280, 21191, 24536, 27609, 25388, 26336, 24396, 26775, 11514, 0, 5821, 5471, 7860, 4281, 4915, 6558, 5395, 5509, 5299, 6497, 1318, 2152, 5535, 3738, 4605, 4057, 4504, 3985, 4852, 2140, 0, 266, 0, 76, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 301, 0, 1097, 0, 7512, 10349, 7680, 17157, 20731, 20823, 17866, 19375, 18926, 18983, 18990, 18337, 17932, 18150, 18433, 20121, 22128, 20898, 21649, 21947, 20112, 20713, 19240, 22693, 25420, 24179, 24780, 24368, 24768, 24213, 25221, 22422, 20291, 12323, 10417, 16117, 16797, 6793, 0, 808, 0, 222, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 266, 0, 901, 0, 7292, 16404, 10411, 9532, 3061, 0, 333, 0, 100, 0, 1, 12, 0, 579, 3188, 3345, 3013, 4316, 6446, 9381, 2366, 2476, 10166, 6420, 1123, 46, 1847, 3623, 4741, 4817, 4994, 3087, 1195, 1408, 399, 0, 34, 0, 11, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 139, 0, 578, 0, 4213, 6953, 7073, 0, 10925, 29291, 27497, 30505, 29671, 29981, 29018, 29269, 28813, 29797, 27399, 35940, 16655, 0, 3612, 938, 3863, 2983, 4082, 3826, 3819, 3908, 3381, 4735, 4832, 3975, 4826, 5298, 4278, 3793, 3937, 3715, 4123, 3374, 4773, 1939, 11412, 21981, 21526, 21747, 24236, 11863, 343, 3829, 2984, 5373, 4990, 5905, 2233, 0, 213, 0, 0, 283, 0, 2525, 5830, 5616, 11457, 5155, 0, 632, 0, 190, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 142, 0, 1656, 951, 10110, 19968, 18014, 15332, 23704, 31568, 27623, 26932, 21899, 18646, 19994, 20518, 21417, 21528, 21757, 21255, 22268, 20146, 27157, 33304, 30704, 26523, 33761, 16065, 0, 6029, 3735, 6255, 3701, 6974, 0, 16898, 32178, 22989, 24782, 21653, 21318, 18871, 17965, 14925, 8906, 6678, 6643, 4879, 1576, 0, 165, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 220, 0, 745, 0, 6599, 18317, 17606, 17449, 11782, 9501, 14771, 18037, 19353, 19555, 21088, 22368, 22564, 22925, 22693, 24015, 25719, 26164, 26197, 26496, 26675, 25367, 23683, 23390, 22487, 24233, 24640, 26125, 25856, 31745, 14293, 0, 6574, 5039, 5609, 5498, 5927, 5360, 4792, 5041, 4818, 5118, 4621, 5580, 2466, 0, 306, 0, 87, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 201, 0, 739, 0, 6289, 7752, 10043, 25571, 29380, 27964, 25182, 23136, 22001, 22963, 23318, 25077, 28278, 30227, 28998, 28219, 29508, 30867, 31478, 31423, 31230, 31723, 30743, 32735, 26568, 23168, 26307, 25041, 26694, 32204, 23471, 8070, 6915, 7042, 6264, 4719, 2746, 1283, 1628, 1246, 387, 0, 38, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 303, 0, 1058, 0, 8665, 20427, 18094, 20105, 19299, 19518, 19531, 20414, 20859, 23993, 24168, 22039, 22384, 22058, 22078, 21939, 22915, 23723, 24363, 23347, 25561, 23895, 25455, 10384, 0, 1804, 11496, 25290, 21153, 24882, 12387, 4633, 5088, 548, 2366, 454, 0, 23, 0, 19, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 71, 0, 127, 0, 3120, 14620, 3123, 8736, 27861, 26540, 26940, 20617, 19423, 20666, 20358, 20788, 20514, 20586, 20632, 21010, 21447, 21598, 21847, 21762, 21614, 21712, 21684, 21135, 20056, 19449, 19770, 19304, 20149, 18562, 21759, 11908, 4748, 4570, 15122, 15759, 4210, 6259, 3188, 4389, 2948, 1357, 54, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 34, 0, 120, 0, 791, 791, 0, 120, 0, 34, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 156, 0, 441, 0, 4605, 13047, 416, 9381, 23311, 19751, 21691, 20611, 21200, 20879, 21086, 20781, 20851, 21069, 21268, 21521, 21502, 21463, 21414, 20808, 19842, 19758, 19531, 19245, 19774, 20196, 22417, 26060, 9373, 0, 2470, 4564, 5722, 6112, 6245, 3193, 2828, 3567, 2308, 1844, 2317, 438, 0, 17, 0, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 140, 0, 542, 0, 4467, 10177, 9820, 5704, 16159, 26542, 22104, 21286, 19370, 20456, 20122, 20834, 20865, 21868, 22682, 22687, 22418, 21763, 21901, 21942, 21823, 21634, 20678, 19560, 19803, 19547, 20109, 20072, 24002, 25830, 26170, 29641, 29740, 30008, 29619, 30295, 29047, 31468, 24898, 24278, 17019, 5217, 9596, 6269, 1721, 0, 144, 0, 27, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 208, 0, 726, 0, 5144, 7295, 0, 428, 0, 449, 0, 1211, 0, 9764, 22779, 19920, 21993, 21525, 22500, 22355, 22727, 22712, 22649, 22462, 22175, 22245, 23415, 24310, 23310, 25596, 26765, 26232, 25788, 23704, 16963, 7635, 6302, 7609, 7176, 6710, 6406, 7174, 5756, 7187, 2159, 2006, 3172, 0, 534, 0, 141, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 67, 0, 367, 0, 2527, 4719, 13051, 4192, 10784, 29093, 24098, 26087, 20160, 17323, 17202, 16831, 18728, 18935, 19739, 20509, 20471, 21245, 20590, 21306, 21444, 21458, 22101, 22409, 23052, 23038, 24725, 25449, 25467, 25105, 25918, 24354, 27546, 16493, 2581, 6881, 5338, 4850, 6118, 4775, 3875, 3289, 3763, 1595, 0, 195, 0, 55, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 177, 0, 626, 0, 5133, 11085, 6938, 10189, 20974, 26192, 24857, 25469, 25169, 25283, 25329, 24758, 22907, 21717, 21796, 21622, 20769, 19538, 18524, 17945, 17132, 18053, 17520, 21334, 23863, 25448, 23968, 28939, 16337, 0, 17037, 29176, 18510, 20774, 21296, 20770, 17421, 8941, 3959, 2282, 166, 27, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 86, 0, 295, 0, 3131, 3702, 137, 346, 0, 79, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 285, 0, 1000, 0, 8638, 21538, 16159, 13261, 21636, 29575, 27952, 27925, 26789, 25580, 23915, 23225, 23805, 24172, 23845, 24263, 24481, 22682, 21847, 22376, 21432, 21471, 22574, 22382, 23591, 23228, 26782, 29437, 27664, 27730, 28779, 30304, 30046, 30513, 29690, 31192, 28428, 33954, 15838, 0, 3759, 3016, 1805, 539, 1535, 0, 247, 0, 65, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 253, 0, 945, 0, 6519, 10420, 13944, 25681, 28057, 32194, 31111, 30982, 31465, 30255, 29709, 29825, 30064, 29389, 30761, 28172, 33372, 16262, 0, 4464, 2037, 3327, 1018, 283, 1589, 3123, 2313, 5910, 0, 15922, 28910, 21228, 24678, 21842, 20743, 17218, 15885, 5692, 0, 1890, 283, 9, 0, 0, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 233, 0, 832, 0, 8584, 15103, 13898, 16241, 15719, 26192, 30702, 30147, 30385, 29296, 28610, 24131, 21064, 22914, 23700, 24064, 24287, 25235, 25568, 26515, 27110, 26742, 22008, 30960, 14769, 0, 4459, 2351, 3381, 3214, 2311, 5740, 0, 16484, 33165, 20601, 21438, 19858, 20597, 19805, 20928, 18981, 22838, 10127, 0, 1327, 0, 609, 0, 2378, 5308, 4453, 1633, 0, 191, 0, 43, 0, 0, 46, 0, 431, 916, 205, 0, 11, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 109, 0, 285, 0, 6813, 14298, 2704, 6514, 16818, 24501, 28628, 25815, 22844, 18460, 20331, 19622, 20177, 20028, 20077, 19546, 20887, 22736, 22753, 22866, 22753, 22907, 22645, 23405, 24383, 26457, 29972, 21105, 5804, 0, 8703, 20494, 17892, 24042, 25245, 19309, 21316, 9423, 73, 2624, 1142, 1863, 1111, 1456, 668, 2039, 1424, 0, 203, 0, 57, 0, 8, 0, 0, 12, 0, 40, 0, 529, 2310, 2902, 2807, 2791, 2903, 2651, 3183, 1411, 0, 175, 0, 50, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 444, 0, 1528, 0, 12570, 29134, 21075, 21415, 20551, 20206, 20400, 20804, 21911, 22864, 22010, 20933, 20173, 20059, 21233, 21651, 22336, 22609, 23121, 22749, 22388, 22728, 26561, 27107, 29304, 24449, 36625, 11837, 12431, 32358, 18405, 15362, 683, 9547, 7855, 3459, 4908, 3653, 3751, 3655, 3626, 3799, 3442, 4155, 1836, 0, 228, 0, 65, 0, 15, 0, 3, 0, 5, 0, 215, 1215, 629, 0, 79, 0, 23, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 169, 0, 609, 0, 5043, 11506, 8686, 9353, 18424, 25092, 20603, 19614, 20746, 20246, 19514, 19842, 20585, 20759, 21399, 21606, 21527, 22525, 23007, 22724, 22561, 22456, 22291, 22326, 22314, 22354, 22236, 22410, 23382, 29925, 13897, 584, 7040, 7111, 6142, 5435, 6679, 5612, 5473, 5626, 5895, 2697, 0, 3110, 2710, 0, 394, 0, 114, 0, 23, 0, 0, 0, 12, 0, 70, 0, 251, 0, 1636, 1768, 504, 1498, 148, 23, 0, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 108, 0, 402, 0, 3263, 8287, 10921, 9534, 6251, 7205, 6987, 6627, 7691, 5334, 13221, 20697, 17091, 17659, 17872, 18035, 18690, 20588, 21601, 22497, 22831, 22892, 22770, 21396, 24754, 27469, 26540, 26170, 25993, 27972, 27355, 28766, 22716, 18932, 18591, 16769, 10491, 2246, 9827, 17831, 6687, 0, 722, 0, 212, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 194, 0, 652, 0, 5627, 14169, 10684, 15431, 20151, 26367, 31605, 31006, 29323, 26233, 25747, 25253, 24053, 21830, 20001, 19160, 17990, 17059, 16860, 17005, 17730, 20941, 20439, 20182, 21522, 23296, 9112, 0, 1192, 0, 402, 113, 7, 836, 763, 0, 114, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 69, 0, 246, 0, 2371, 6117, 3086, 5315, 20523, 29512, 28601, 28644, 28370, 28769, 28794, 28743, 29059, 28334, 29728, 27135, 32319, 15339, 0, 4410, 2687, 4694, 3774, 4118, 4432, 4055, 4762, 5849, 5067, 4224, 4450, 5807, 2915, 5979, 0, 16849, 28077, 13592, 12872, 11895, 20924, 21528, 22641, 22497, 24155, 12068, 1363, 4509, 2081, 2996, 1196, 0, 149, 0, 49, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 107, 0, 919, 2625, 4899, 6479, 11027, 15231, 10757, 16384, 17393, 22640, 32650, 31597, 29999, 26910, 28129, 29184, 27051, 29538, 28389, 35848, 16677, 0, 2945, 270, 2264, 1849, 1462, 407, 1449, 3044, 5192, 5580, 6206, 4413, 6772, 0, 17345, 31507, 20871, 23916, 21883, 23331, 21930, 24025, 17697, 10649, 8591, 5628, 2663, 0, 343, 0, 68, 0, 11, 0, 0, 2, 0, 7, 0, 48, 48, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 48, 804, 9684, 17132, 14771, 12681, 12771, 17938, 19731, 19390, 20965, 20918, 22283, 23279, 22395, 22876, 24569, 24889, 25048, 24984, 25024, 24979, 25066, 24825, 24789, 23722, 25860, 25196, 28073, 25582, 28123, 22475, 4738, 6023, 6671, 5903, 5880, 5371, 6253, 2786, 0, 276, 0, 80, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 91, 0, 311, 0, 4518, 21651, 29986, 27232, 26287, 23426, 21601, 22474, 23258, 24759, 26650, 29201, 28551, 28183, 28551, 29274, 30618, 32194, 28870, 24254, 23381, 22823, 22908, 23958, 24346, 25773, 26804, 26395, 28795, 33680, 26341, 10955, 7256, 6709, 4229, 2396, 1626, 1422, 1405, 1423, 1393, 1463, 1329, 1601, 708, 0, 88, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 79, 0, 193, 0, 2924, 14305, 14056, 14012, 2957, 8019, 23883, 18971, 20401, 19822, 20120, 20267, 20059, 20218, 20811, 23727, 26347, 26377, 25262, 23965, 24027, 24174, 24087, 24217, 23997, 24347, 23724, 25495, 22633, 6170, 799, 3523, 13745, 24682, 16423, 6988, 4821, 3060, 1240, 1833, 630, 0, 57, 0, 20, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 0, 60, 0, 413, 773, 1408, 826, 0, 113, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 227, 0, 795, 0, 6275, 13471, 10596, 11832, 11356, 11262, 11958, 10276, 15980, 21507, 19759, 20802, 21016, 21713, 21624, 22592, 23379, 23601, 23739, 22742, 22865, 22989, 22303, 22693, 21962, 22145, 21276, 23456, 25652, 27495, 15101, 5703, 9570, 7052, 6936, 7094, 6448, 5308, 4753, 4200, 3671, 1571, 54, 26, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 21, 0, 76, 0, 503, 503, 0, 76, 0, 21, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 157, 0, 448, 0, 4699, 13419, 716, 9243, 24830, 22401, 21476, 18851, 20266, 20151, 20048, 19616, 20129, 21983, 22394, 22076, 22625, 22831, 22464, 22018, 22242, 21769, 21172, 21287, 21222, 21467, 21834, 21887, 22047, 21666, 22409, 21025, 23809, 14420, 3114, 3945, 1652, 1924, 1048, 1937, 2709, 730, 0, 60, 0, 20, 0, 5, 0, 0, 0, 0, 8, 0, 49, 0, 179, 0, 2482, 6059, 7751, 8517, 7963, 5759, 1133, 0, 74, 0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 0, 88, 0, 1656, 8902, 14112, 1047, 9360, 25781, 19403, 19148, 20036, 20332, 20259, 20315, 20199, 20451, 19900, 21727, 23545, 23047, 23339, 23535, 23585, 23510, 23609, 22828, 22595, 22597, 22585, 23567, 26831, 28001, 29582, 25642, 21217, 10095, 938, 6448, 7049, 7592, 11526, 16920, 17785, 16577, 20966, 10799, 0, 540, 0, 169, 0, 29, 0, 0, 0, 17, 0, 85, 0, 301, 0, 2340, 4790, 3198, 1306, 0, 167, 0, 42, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29729, 28756, 29021, 29343, 30109, 29864, 29423, 27373, 27753, 17661, 9426, 11332, 9064, 6439, 4361, 4827, 3119, 6387, 7639, 6223, 6971, 6350, 6710, 6393, 6799, 6141, 7409, 3277, 0, 407, 0, 116, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 154, 0, 533, 0, 4646, 12324, 11273, 11319, 11286, 11074, 11622, 10547, 12711, 5620, 0, 698, 0, 199, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 199, 200, 0, 32, 0, 0, 120, 0, 460, 0, 1583, 0, 12871, 29604, 30924, 29377, 37992, 12439, 11661, 38288, 26198, 29305, 27240, 27839, 26824, 27092, 27547, 27691, 27848, 27791, 27466, 26958, 27007, 27175, 27125, 26867, 27139, 27334, 27275, 27427, 27171, 27349, 27232, 27054, 27219, 27327, 27337, 27250, 27077, 26895, 26884, 26871, 26897, 26849, 26936, 26761, 27369, 28269, 28450, 28514, 28168, 28312, 28849, 28833, 28558, 27444, 25123, 9013, 0, 718, 0, 164, 0, 0, 264, 0, 3131, 8342, 8559, 11200, 6975, 5279, 3148, 0, 458, 0, 123, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 449, 634, 1453, 3341, 8059, 11616, 11241, 12403, 12264, 12519, 13705, 12100, 9592, 8656, 8837, 8839, 8689, 9062, 8007, 8427, 9288, 9248, 6665, 1094, 0, 43, 0, 17, 0, 10, 0, 17, 0, 182, 572, 215, 0, 42, 0, 102, 0, 348, 0, 2802, 6309, 5676, 5441, 8896, 17607, 22605, 24389, 24662, 24549, 24327, 24527, 24536, 24866, 25144, 25219, 24849, 25715, 23906, 28525, 28250, 34547, 17061, 0, 4842, 0, 15828, 33760, 28054, 29080, 26896, 29104, 28852, 29727, 29780, 30184, 29896, 29055, 28604, 27906, 26215, 25357, 24622, 24492, 22413, 20564, 20555, 20388, 21069, 22742, 23853, 23174, 22578, 21262, 18240, 15194, 5986, 317, 1920, 1104, 1598, 1240, 1620, 688, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 97, 0, 788, 1770, 1488, 1597, 1597, 1488, 1770, 763, 0, 0, 180, 0, 815, 0, 7184, 19632, 23131, 28363, 30291, 31653, 31480, 31327, 31073, 30188, 28701, 28755, 29537, 30297, 29666, 24109, 6843, 0, 652, 0, 126, 0, 0, 387, 0, 3492, 10080, 17192, 25593, 26916, 28239, 28799, 28649, 28748, 28657, 28757, 28596, 29041, 29288, 29100, 29251, 28884, 29315, 27386, 30344, 24922, 36642, 12715, 11229, 35291, 26052, 25004, 17195, 20176, 18045, 17535, 17110, 16819, 16744, 15639, 13810, 13981, 12987, 12027, 11634, 13314, 17201, 20289, 18056, 10091, 0, 21398, 20210, 0, 3028, 0, 862, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 98, 0, 860, 3663, 12413, 19618, 21657, 23747, 25181, 29501, 26490, 34020, 15395, 0, 3124, 474, 2480, 1666, 2125, 2079, 1655, 2143, 177, 2689, 0, 14922, 33484, 27753, 30665, 28562, 28927, 28694, 28846, 28728, 29147, 29912, 29825, 29906, 29877, 30477, 30977, 30853, 30866, 30947, 30742, 31186, 29700, 28311, 29043, 28972, 28897, 29420, 28322, 27350, 27860, 27950, 28367, 28566, 28565, 29118, 29502, 29510, 29114, 26687, 25628, 23871, 22411, 18998, 15932, 17227, 13943, 3746, 0, 365, 0, 206, 0, 1000, 2973, 5729, 6937, 8708, 6826, 4477, 5936, 5318, 5624, 5492, 5502, 5634, 4718, 1237, 0, 110, 0, 32, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 63, 0, 217, 0, 3282, 16384, 24411, 26399, 27429, 27619, 28452, 28576, 28789, 28482, 29244, 28456, 30417, 26234, 35154, 11226, 11131, 35139, 26550, 30665, 27823, 28655, 28226, 28069, 28043, 27924, 27671, 27087, 26727, 26555, 25993, 25995, 25918, 25756, 25848, 25735, 25911, 25583, 26667, 27935, 27699, 28624, 28757, 29185, 29460, 29372, 29122, 28990, 29295, 29199, 29462, 28562, 28209, 28308, 28284, 28496, 27945, 26225, 25554, 25371, 24331, 19696, 19266, 7730, 0, 935, 0, 311, 0, 219, 0, 1337, 2965, 2562, 3140, 3477, 3217, 2823, 2880, 2964, 2720, 3257, 1446, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 181, 0, 644, 0, 5590, 15414, 18416, 21927, 22115, 23000, 24139, 24678, 26925, 28990, 29354, 30287, 30529, 31270, 32736, 30316, 28103, 28985, 28669, 28927, 28812, 28898, 29066, 29242, 29244, 29119, 29017, 29002, 29109, 29060, 29175, 29091, 29070, 29080, 29416, 29604, 29615, 29759, 29691, 29741, 29677, 29798, 29551, 30079, 28237, 22424, 6732, 0, 688, 0, 195, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 105, 0, 370, 0, 2940, 6755, 6916, 9300, 8598, 10484, 11568, 10073, 10178, 8487, 6650, 7166, 4528, 2479, 3100, 2730, 3041, 2677, 3275, 1438, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 294, 0, 1019, 0, 8470, 19456, 15891, 19699, 27043, 26961, 34882, 17080, 0, 4858, 0, 16487, 33604, 27260, 30332, 28353, 29267, 28868, 29213, 29250, 29259, 29179, 28921, 29078, 29193, 29152, 29192, 29134, 29232, 29046, 29598, 29849, 29653, 29836, 29886, 29789, 29651, 30125, 29869, 29617, 28734, 27427, 24015, 25256, 14999, 773, 261, 0, 92, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 86, 0, 310, 0, 2330, 4340, 3446, 3700, 3914, 1910, 0, 246, 0, 66, 0, 0, 63, 0, 353, 0, 1250, 0, 9978, 22754, 22543, 27475, 26185, 26737, 26772, 27588, 27786, 27843, 27737, 27664, 27731, 28081, 28284, 28306, 27896, 27048, 26932, 25972, 25259, 25477, 25342, 25465, 25298, 25601, 24666, 23170, 20579, 22430, 26477, 27644, 28501, 28471, 28440, 28706, 28207, 29436, 26860, 32802, 14354, 0, 3843, 1917, 2013, 4528, 0, 16727, 36685, 30362, 32253, 29576, 30273, 29576, 28382, 23000, 19920, 17664, 12005, 10252, 10627, 10158, 9609, 9073, 9185, 8922, 9402, 8527, 10275, 4546, 0, 564, 0, 161, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 134, 0, 521, 0, 7059, 23692, 28677, 30816, 29245, 36487, 16512, 0, 4430, 1399, 3171, 2226, 2136, 1707, 1881, 1879, 2312, 2663, 2873, 2916, 3086, 3002, 3038, 3088, 2942, 2827, 2961, 3092, 2779, 2965, 2902, 3214, 4256, 4613, 4466, 4717, 4184, 5250, 3232, 7135, 0, 14695, 32988, 26711, 30097, 28528, 29147, 28531, 28844, 29161, 29286, 28761, 30004, 28750, 28815, 19800, 3371, 0, 149, 0, 47, 0, 5, 0, 0, 68, 0, 239, 0, 2139, 6099, 7060, 7983, 8212, 8006, 8398, 8053, 7153, 7533, 7188, 7647, 6899, 8333, 3683, 0, 457, 0, 130, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2607, 2603, 2628, 2569, 2733, 2595, 2206, 2342, 2401, 1956, 1903, 2367, 2721, 2677, 2807, 2675, 2664, 1122, 0, 264, 0, 1111, 2469, 2648, 2983, 3133, 1637, 0, 1595, 1326, 0, 191, 0, 59, 0, 27, 0, 52, 0, 462, 1199, 809, 613, 705, 575, 799, 362, 1792, 3362, 3154, 3294, 2794, 2730, 2959, 2728, 3167, 3662, 3459, 3569, 3536, 3573, 3634, 3644, 3658, 3579, 3514, 3486, 3554, 3510, 3727, 3335, 3145, 1245, 0, 149, 0, 42, 0, 8, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1285, 2965, 2562, 2868, 2825, 3209, 3370, 3459, 3301, 3306, 2863, 2350, 2397, 2337, 2322, 2327, 2576, 2591, 2584, 2690, 2645, 3075, 3563, 3646, 3751, 3739, 3663, 3749, 3920, 3879, 3913, 4017, 3943, 3919, 3406, 3743, 1539, 0, 185, 0, 57, 0, 33, 0, 77, 0, 699, 2015, 2095, 2642, 2848, 2892, 2953, 3145, 3297, 3609, 3911, 3813, 3824, 3669, 3908, 3479, 2772, 2703, 2764, 2793, 2432, 3042, 3115, 2604, 2838, 2847, 3127, 2943, 3608, 4324, 3625, 3641, 3807, 3733, 3743, 3834, 3976, 3925, 3959, 3927, 3967, 3907, 4008, 3547, 2777, 3064, 994, 0, 0, 1423, 3447, 2926, 3416, 3358, 3478, 3283, 3430, 3599, 3668, 3843, 3766, 3720, 3149, 2812, 2975, 2935, 2870, 2950, 2861, 2872, 3102, 3003, 2992, 2901, 2927, 2895, 2841, 2861, 2850, 2955, 2962, 2955, 2976, 2933, 3015, 2850, 3389, 3918, 3746, 3861, 3996, 3990, 3979, 3832, 3529, 3766, 3722, 3507, 3274, 3164, 3274, 3391, 3493, 3466, 3450, 3387, 3551, 3630, 3747, 3890, 4122, 3965, 3821, 3441, 2928, 2930, 2705, 2616, 2702, 2742, 2715, 2850, 2728, 2730, 2849, 2807, 2829, 2818, 2822, 2823, 2826, 2891, 2891, 3252, 3685, 3601, 3812, 4042, 3996, 4113, 4198, 4253, 4290, 4082, 4147, 4156, 3827, 4136, 3845, 3307, 3282, 3287, 3437, 3434, 3410, 3289, 3320, 3279, 3532, 3670, 3673, 3894, 3721, 3713, 3101, 2719, 2902, 2689, 2656, 2650, 2661, 2643, 2677, 2608, 2838, 3095, 3111, 3125, 2975, 2869, 2700, 2676, 2797, 2596, 2995, 3471, 3481, 3466, 3472, 3755, 3746, 4134, 4552, 4617, 4603, 4528, 4531, 4538, 4169, 3749, 3590, 3277, 3268, 3285, 3134, 3157, 3377, 3340, 3264, 3413, 3301, 3450, 3619, 3576, 3581, 3610, 3536, 3695, 3165, 2649, 2928, 2952, 3180, 3119, 3111, 3174, 2888, 2862, 2932, 2823, 2864, 2804, 3206, 3626, 3560, 3600, 3713, 3672, 3748, 3837, 4291, 4683, 4653, 4774, 4883, 4740, 4700, 4885, 5380, 2045, 0, 290, 0, 756, 2622, 2718, 2278, 2407, 2365, 2350, 2431, 2234, 2895, 3500, 3467, 3446, 3447, 3647, 3593, 3175, 2997, 3301, 3184, 3157, 3320, 3198, 2691, 2536, 2610, 2418, 2361, 2750, 2747, 3149, 3461, 3451, 3564, 3548, 3800, 4020, 4158, 4504, 4849, 4687, 4894, 4166, 3446, 3532, 3541, 3850, 3828, 3897, 3775, 3999, 3583, 4412, 1830, 41, 598, 0, 0, 947, 2332, 1968, 2535, 2698, 2807, 2958, 3171, 3322, 3199, 3096, 3198, 2794, 2611, 2813, 2776, 2347, 1898, 1901, 2134, 2126, 2084, 2933, 2866, 2888, 3471, 3461, 3613, 3825, 4131, 4195, 4327, 3985, 3692, 3772, 3744, 3738, 3781, 3682, 4025, 4386, 3910, 4106, 3937, 4670, 1999, 0, 239, 0, 361, 808, 205, 482, 1898, 1875, 2311, 2894, 2946, 3043, 3215, 3393, 3523, 3572, 3459, 3339, 2995, 3055, 1274, 0, 767, 1422, 1478, 1894, 2663, 3082, 3007, 3337, 3503, 3459, 3485, 3461, 3492, 3440, 3573, 3593, 3728, 4011, 4047, 4270, 4041, 3832, 4474, 4037, 4667, 2051, 0, 255, 0, 73, 0, 14, 0, 3, 0, 13, 0, 219, 1263, 2507, 2984, 3053, 3159, 3215, 3334, 3269, 3369, 3078, 2862, 1212, 0, 907, 1695, 1482, 1623, 1477, 1681, 1317, 2487, 3844, 3758, 3918, 3700, 3683, 3446, 3580, 3842, 3840, 3897, 4077, 3828, 3718, 4283, 4141, 4540, 1782, 0, 210, 0, 60, 0, 11, 0, 0, 7, 0, 30, 0, 239, 707, 1827, 2918, 3003, 3113, 3176, 3358, 3414, 3410, 3395, 3432, 3355, 3514, 2998, 2459, 2374, 2762, 3302, 3082, 3322, 3634, 3645, 3789, 3856, 3449, 3671, 3451, 3731, 4101, 3861, 4196, 4136, 4151, 4298, 3821, 3647, 1364, 0, 158, 0, 45, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 57, 0, 198, 0, 1686, 4066, 2623, 1909, 2272, 1094, 0, 958, 2602, 805, 467, 2357, 2648, 2860, 3129, 3519, 3621, 3925, 3868, 3623, 1226, 0, 134, 0, 38, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 43, 0, 151, 0, 1261, 3067, 2818, 3081, 3277, 3727, 3720, 3753, 3682, 3550, 2851, 2622, 3014, 2730, 2714, 2732, 2528, 1975, 1991, 2294, 2362, 2488, 2958, 3456, 3499, 3642, 3758, 3739, 3526, 1189, 0, 129, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1309, 3083, 2367, 2857, 3328, 3503, 3485, 3527, 3674, 2519, 2170, 2806, 2438, 2502, 2931, 2804, 2836, 2952, 2985, 2783, 2548, 2848, 2134, 2085, 2400, 2392, 2706, 2688, 3101, 3333, 3467, 3700, 3724, 3817, 3699, 3902, 3536, 4262, 1885, 0, 234, 0, 62, 0, 0, 38, 0, 157, 0, 1291, 3082, 2892, 3351, 3233, 3409, 3391, 3439, 3183, 2353, 2047, 2147, 2106, 2471, 2617, 2601, 2867, 2904, 2945, 2904, 2999, 2993, 3037, 3100, 3113, 3177, 3157, 3190, 3172, 3191, 3163, 3217, 3105, 3458, 3711, 3875, 3631, 4087, 1743, 0, 213, 0, 60, 0, 23, 0, 55, 0, 198, 0, 1535, 3184, 2688, 3264, 3338, 3279, 3075, 3388, 3417, 806, 746, 2671, 2388, 2739, 2891, 3131, 3090, 3141, 3205, 3202, 3278, 3305, 3300, 3291, 3317, 3263, 3372, 3062, 2957, 2587, 2304, 2554, 2654, 2655, 3131, 3661, 3410, 3606, 3396, 3877, 1569, 0, 187, 0, 60, 0, 42, 0, 112, 0, 928, 2347, 2663, 3253, 3125, 3577, 3298, 3287, 3174, 2680, 2426, 2160, 2705, 2798, 2667, 2680, 2664, 2679, 2664, 2684, 2646, 2802, 3136, 2995, 2962, 3050, 3042, 3091, 2938, 2810, 2708, 2718, 2749, 2786, 2771, 2844, 2873, 3252, 3614, 3516, 3579, 3429, 3444, 2867, 2792, 1143, 0, 112, 0, 0, 155, 0, 1446, 3469, 3085, 3451, 3339, 3584, 3369, 3097, 3229, 3077, 3308, 2915, 3660, 1402, 435, 2659, 369, 867, 2333, 1965, 2349, 2473, 2462, 2161, 1735, 2102, 883, 0, 66, 15, 0, 698, 2162, 2158, 2713, 3194, 3264, 3542, 3490, 3727, 3390, 2665, 894, 0, 99, 0, 27, 0, 5, 0, 0, 9, 0, 39, 0, 120, 0, 1186, 3394, 1121, 0, 0, 445, 1575, 1813, 2313, 2622, 2539, 2648, 2853, 2764, 2505, 2510, 2230, 2159, 868, 0, 93, 0, 0, 276, 1447, 1971, 2544, 3068, 3161, 3364, 3536, 3491, 3645, 3341, 4500, 2102, 0, 265, 0, 76, 0, 12, 0, 0, 18, 0, 65, 0, 656, 2240, 2733, 2464, 2465, 2800, 2468, 2351, 768, 0, 0, 742, 2480, 2472, 2438, 2234, 2817, 1208, 0, 153, 0, 66, 0, 92, 0, 725, 1943, 2097, 2604, 3124, 3496, 3423, 3426, 3580, 3619, 3653, 3560, 3745, 3398, 4093, 1811, 0, 225, 0, 64, 0, 10, 0, 0, 35, 0, 133, 0, 857, 967, 1037, 2248, 2152, 2532, 2135, 2653, 1100, 0, 90, 10, 0, 536, 564, 0, 76, 0, 0, 34, 0, 405, 1063, 901, 1713, 2244, 2092, 2178, 2112, 2181, 2077, 2454, 3322, 3426, 3569, 3555, 4068, 1647, 0, 196, 0, 56, 0, 11, 0, 0, 0, 0, 0, 0, 0, 3, 0, 8, 0, 15, 0, 424, 2216, 1116, 0, 140, 0, 41, 0, 9, 0, 0, 0, 10, 0, 47, 0, 160, 0, 1413, 3532, 2204, 2589, 4061, 3174, 3091, 3816, 3322, 3472, 3740, 3682, 3620, 2885, 3672, 1737, 0, 221, 0, 63, 0, 12, 0, 0, 0, 3, 0, 13, 0, 46, 0, 427, 1188, 1080, 1652, 2702, 2678, 2118, 2012, 2045, 1989, 2092, 1903, 2278, 1029, 0, 187, 0, 673, 2148, 2633, 2571, 3284, 1190, 0, 0, 1661, 3948, 3076, 3473, 3550, 3427, 3819, 1552, 0, 184, 0, 53, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 93, 0, 787, 2019, 1704, 2587, 1112, 0, 79, 31, 0, 1002, 3045, 2246, 1954, 821, 0, 104, 0, 30, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 0, 42, 0, 554, 2079, 890, 0, 103, 0, 31, 0, 7, 0, 0, 6, 0, 24, 0, 74, 0, 778, 2400, 889, 0, 94, 0, 29, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 55, 0, 895, 1603, 389, 0, 27, 0, 9, 0, 3, 0, 0, 0, 0, 0, 2, 0, 5, 0, 12, 0, 288, 1449, 718, 0, 89, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 25, 0, 90, 0, 595, 595, 0, 90, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 198, 198, 0, 30, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 19, 0, 68, 0, 450, 450, 0, 68, 0, 19, 0, 3, 0, 0, 0, 0, 0, 1, 0, 5, 0, 19, 0, 125, 125, 0, 19, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 633, 1429, 2018, 2193, 2176, 2138, 2240, 2037, 2451, 1085, 0, 134, 0, 38, 0, 7, 0, 1, 0, 8, 0, 28, 0, 424, 321, 0, 46, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 44, 0, 147, 0, 1224, 2670, 631, 0, 40, 0, 15, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 47, 0, 175, 0, 1129, 962, 39, 1004, 2360, 3010, 2596, 2805, 692, 0, 56, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 60, 0, 218, 0, 1457, 1475, 0, 599, 1961, 1133, 0, 147, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 56, 0, 206, 0, 1345, 1250, 0, 0, 651, 815, 0, 126, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1545, 1610, 1540, 1582, 1739, 1395, 2115, 740, 3287, 0, 14847, 31206, 25333, 28322, 26995, 26416, 27153, 24572, 24692, 10264, 0, 1048, 0, 301, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 86, 338, 214, 277, 251, 66, 132, 97, 117, 104, 115, 85, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 883, 0, 3138, 0, 20590, 20829, 0, 4379, 0, 2528, 1622, 2417, 2410, 2739, 3011, 3195, 2770, 2929, 3393, 3468, 3258, 3103, 3078, 2897, 2915, 2764, 2726, 2823, 2505, 2027, 1547, 1459, 1358, 1269, 1416, 1452, 1526, 1480, 1541, 1439, 1621, 1260, 2459, 3790, 3566, 3594, 3562, 3830, 3453, 3247, 3190, 3149, 3104, 2694, 2150, 634, 0, 64, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 30, 551, 1092, 1456, 1663, 1623, 1676, 1587, 1798, 1898, 1799, 1453, 1957, 644, 2210, 281, 7254, 16774, 15160, 17118, 19362, 21795, 22140, 21917, 23356, 24622, 23248, 22432, 23053, 20738, 24381, 10669, 0, 1983, 110, 1082, 639, 960, 827, 847, 901, 786, 1003, 566, 2021, 3544, 2950, 3484, 3801, 4065, 4148, 4260, 4227, 4182, 4219, 4130, 3927, 3861, 4049, 3818, 3635, 3543, 3330, 2873, 2184, 1656, 523, 0, 55, 0, 15, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 276, 0, 984, 0, 9449, 20790, 21221, 23631, 23583, 25941, 25032, 25743, 25783, 26446, 26853, 27422, 27371, 26713, 27220, 26444, 27800, 25349, 30207, 14310, 0, 3117, 688, 3432, 3786, 4028, 4341, 4403, 4496, 4355, 4151, 4178, 4107, 4127, 4211, 4169, 4263, 4387, 4188, 4417, 4298, 4450, 4557, 4314, 4482, 4498, 4532, 4234, 4150, 4002, 4104, 3705, 3688, 1507, 0, 182, 0, 51, 0, 10, 0, 39, 0, 195, 0, 689, 0, 5565, 13113, 11388, 12682, 12055, 14342, 5546, 0, 653, 0, 193, 0, 54, 0, 170, 708, 1011, 1091, 1075, 1203, 1281, 1410, 1079, 748, 312, 0, 39, 0, 10, 0, 1, 0, 0, 0, 12, 0, 62, 0, 219, 0, 1793, 4282, 4181, 4679, 4501, 4836, 4906, 4797, 4794, 4585, 4060, 4436, 3718, 2846, 3159, 2734, 3377, 4525, 4663, 4997, 4950, 4613, 4682, 4317, 2410, 1258, 1442, 1348, 1429, 1537, 1480, 1593, 1682, 1813, 1768, 2458, 4236, 4767, 4660, 4700, 4689, 4676, 4727, 4500, 4064, 4164, 4071, 3771, 3344, 2968, 1763, 235, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 887, 0, 3151, 0, 20641, 20627, 0, 3857, 0, 1822, 533, 1124, 253, 0, 6, 32, 0, 245, 0, 884, 0, 7520, 19357, 20143, 22759, 24573, 26205, 26960, 26828, 27012, 23850, 25824, 11483, 0, 2509, 575, 1731, 1088, 1475, 1381, 1997, 2724, 3258, 3551, 3733, 4461, 4767, 4837, 4876, 5043, 5114, 5163, 5199, 5152, 5240, 5287, 5497, 5608, 5570, 5602, 5560, 5636, 5358, 4787, 4646, 4606, 4628, 4438, 4300, 3912, 3562, 1260, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 194, 0, 910, 0, 7333, 23432, 30566, 29528, 36790, 16379, 0, 2887, 314, 2322, 1942, 2069, 1527, 1895, 1077, 1916, 340, 2954, 0, 16469, 36143, 29004, 33121, 29262, 30892, 13262, 0, 3764, 2046, 3193, 2549, 2995, 3007, 3056, 3059, 3053, 3062, 3045, 3080, 2953, 2727, 2643, 2935, 3263, 3515, 3853, 4038, 4192, 4104, 4018, 4104, 4195, 3986, 3609, 1193, 0, 128, 0, 37, 0, 0, 47, 0, 252, 0, 875, 0, 7329, 17960, 15543, 16260, 15845, 15557, 15066, 15214, 15368, 14658, 13946, 14314, 13849, 14609, 13266, 15907, 7366, 0, 2657, 1697, 2230, 1674, 1894, 1771, 2020, 2169, 919, 304, 687, 112, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 4, 0, 137, 880, 1452, 1891, 2471, 2694, 2803, 2933, 3151, 3227, 3192, 3202, 3205, 3188, 3226, 3147, 3385, 3547, 3791, 4009, 3985, 4399, 4453, 3806, 3213, 3444, 3379, 3379, 2237, 975, 892, 1090, 1345, 2080, 3193, 3645, 4219, 4647, 4602, 4556, 4821, 4842, 4778, 4832, 4915, 4977, 4872, 4726, 4708, 4767, 4695, 4500, 4626, 4113, 3682, 3819, 3733, 3813, 3708, 3894, 3292, 2529, 2209, 1746, 606, 0, 67, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 92, 220, 163, 224, 131, 291, 0, 1010, 2165, 2044, 2029, 1710, 1740, 1977, 2078, 2117, 2026, 1882, 2068, 2401, 2544, 2596, 2576, 2599, 2541, 2431, 2662, 2388, 2322, 1976, 1620, 1690, 548, 0, 87, 0, 339, 1126, 1710, 2197, 2538, 2856, 3037, 3215, 3267, 3216, 3271, 3176, 3347, 3034, 3657, 1617, 0, 200, 0, 57, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 100, 0, 943, 2434, 2806, 3212, 3539, 2237, 857, 0, 1387, 0, 9904, 25243, 26922, 29474, 28436, 29034, 28601, 29074, 28318, 30618, 32815, 31923, 32079, 30119, 28452, 10519, 0, 2347, 581, 2176, 3275, 4210, 4440, 4368, 4328, 4374, 4241, 4064, 4087, 4226, 4334, 4421, 4479, 4502, 4366, 3977, 4012, 4185, 4151, 4153, 4165, 4164, 4036, 3890, 3804, 3724, 3657, 3632, 3678, 3580, 3769, 3419, 4119, 1822, 0, 226, 0, 64, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 13, 0, 44, 0, 465, 1638, 1914, 1984, 2163, 2288, 2618, 2560, 2696, 3017, 2815, 2858, 3051, 3084, 2901, 2907, 2822, 2751, 2778, 2715, 2941, 3138, 3166, 3163, 3166, 3161, 3172, 3145, 3254, 3367, 2820, 1793, 1342, 476, 0, 54, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 5, 1, 348, 1292, 584, 880, 0, 14875, 26450, 28530, 29079, 35789, 16866, 0, 3612, 541, 2147, 1040, 2028, 981, 1755, 0, 2375, 0, 16422, 36997, 30212, 33790, 27587, 30916, 13334, 0, 2196, 0, 1112, 295, 868, 243, 1921, 3709, 3310, 3494, 3393, 3664, 3595, 3606, 3785, 3733, 3655, 3610, 3519, 3375, 3378, 3335, 3092, 2921, 2241, 1865, 713, 0, 84, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 320, 0, 1113, 0, 8993, 20381, 16893, 18804, 15448, 4733, 0, 474, 0, 130, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 307, 0, 1061, 0, 9357, 25538, 25071, 28260, 29472, 30450, 31537, 31538, 31427, 31296, 31309, 31326, 31316, 31317, 30782, 27769, 28017, 11117, 0, 2517, 613, 2176, 2609, 3051, 3338, 2988, 2789, 2857, 2570, 2643, 2817, 2884, 2997, 3076, 3228, 3276, 3363, 3520, 3665, 3598, 3506, 3413, 3277, 2570, 1996, 2054, 653, 0, 66, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 0, 528, 0, 1857, 0, 14949, 34024, 29594, 32311, 30364, 30439, 28447, 28238, 27533, 28158, 27521, 25961, 8989, 0, 947, 0, 273, 0, 56, 0, 0, 0, 3, 0, 12, 0, 100, 91, 0, 13, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 382, 0, 1348, 0, 10818, 25212, 22403, 25700, 23018, 24812, 9333, 0, 1094, 0, 315, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 594, 1147, 1324, 1383, 1752, 1969, 1662, 1643, 1515, 1376, 1736, 1728, 1578, 1807, 1896, 1977, 1888, 1740, 1821, 2125, 2073, 2199, 1577, 1247, 646, 0, 88, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 170, 0, 884, 0, 3139, 0, 20588, 20803, 0, 4283, 0, 899, 0, 156, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 0, 381, 0, 1335, 0, 11405, 29672, 29548, 31572, 30832, 32072, 31696, 31622, 31520, 31059, 30098, 28744, 27053, 25534, 9092, 0, 1671, 318, 1245, 1003, 2198, 3164, 3449, 3575, 3783, 3898, 3722, 3728, 3747, 3678, 3589, 3544, 3596, 3497, 3683, 3340, 4024, 1780, 0, 221, 0, 63, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 189, 0, 668, 0, 7176, 19797, 24363, 28340, 28320, 29325, 29095, 29193, 29219, 29074, 28868, 29107, 24437, 26692, 11632, 0, 1373, 0, 391, 0, 92, 0, 1, 0, 7, 0, 173, 996, 1382, 1268, 1354, 1250, 1410, 1113, 2061, 2974, 2697, 2961, 2809, 2846, 2778, 2664, 2663, 2625, 2367, 1471, 317, 0, 24, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 137, 892, 1267, 1409, 576, 0, 70, 0, 21, 0, 15, 31, 97, 76, 174, 289, 252, 272, 259, 271, 253, 310, 378, 342, 219, 221, 31, 481, 1351, 1760, 1787, 1525, 1551, 1608, 1928, 2037, 1828, 615, 0, 67, 0, 19, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28246, 28894, 29871, 29592, 29574, 29422, 29624, 27441, 27776, 20452, 13905, 15694, 15118, 14862, 16180, 10997, 5185, 6593, 6244, 5719, 4473, 4768, 4249, 3637, 1201, 0, 131, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 27, 0, 76, 0, 1045, 4082, 1791, 0, 210, 0, 64, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 27, 0, 236, 563, 167, 36, 0, 249, 0, 2575, 2065, 8893, 14152, 10732, 14941, 19266, 35918, 15401, 0, 0, 15068, 35811, 26264, 28102, 27291, 28438, 27744, 27343, 27792, 28040, 27600, 27876, 28106, 28191, 28051, 27923, 27661, 27250, 27296, 27494, 27518, 27515, 27523, 27503, 27545, 27462, 27692, 27720, 27756, 27829, 27679, 28034, 27380, 26856, 26947, 27029, 26350, 25574, 25801, 25524, 25074, 25217, 25264, 25477, 25112, 25887, 26912, 26924, 26964, 27742, 24910, 21806, 17309, 4172, 0, 141, 172, 0, 3568, 10602, 7899, 5391, 4665, 4521, 4922, 4815, 4774, 4976, 4532, 5453, 2414, 0, 299, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 175, 0, 603, 0, 5070, 12533, 10668, 11707, 10221, 8437, 8115, 6743, 4447, 3923, 3635, 3306, 3698, 3089, 4229, 1892, 0, 235, 0, 18, 124, 0, 828, 0, 3096, 0, 20038, 18344, 0, 0, 15591, 34302, 15989, 5663, 0, 2112, 0, 7361, 13744, 11780, 13012, 11897, 13315, 10895, 18454, 25809, 22714, 23684, 23777, 23952, 24757, 26195, 28344, 31317, 31123, 33057, 30236, 35857, 16787, 0, 4841, 0, 17460, 35506, 29324, 31337, 28965, 25574, 21656, 22461, 21893, 21412, 21213, 21221, 20966, 20315, 20761, 20786, 21510, 23620, 24270, 24441, 24252, 24349, 24250, 24424, 24089, 24764, 22997, 23134, 19941, 18097, 9821, 0, 500, 0, 144, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 77, 0, 274, 0, 1797, 1797, 0, 272, 0, 59, 0, 0, 139, 0, 893, 1814, 9215, 14822, 15087, 14131, 20620, 26071, 34214, 16688, 0, 5196, 2413, 4078, 3184, 3632, 3560, 3889, 3453, 4090, 2083, 5105, 0, 15741, 34314, 28587, 31467, 29899, 30801, 30170, 30886, 29484, 31361, 29775, 36313, 16115, 0, 2925, 0, 3298, 0, 16933, 36975, 28690, 31133, 27863, 36511, 15848, 0, 2600, 3078, 0, 16450, 36058, 27969, 30646, 25419, 20450, 17715, 16860, 16548, 15798, 15196, 15038, 14298, 12844, 12443, 12022, 11735, 11946, 11602, 12217, 11101, 13319, 6038, 0, 694, 0, 199, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 215, 0, 814, 0, 6711, 15926, 20215, 24401, 33673, 15273, 0, 5040, 2720, 4848, 4207, 4772, 4673, 4918, 4930, 4920, 4592, 5241, 3730, 5877, 397, 16740, 33251, 28153, 30801, 29572, 30213, 29961, 29958, 30186, 29286, 28206, 28281, 28102, 28048, 28005, 27869, 27679, 27852, 27967, 28085, 28408, 28714, 28502, 28486, 28804, 29026, 29185, 29508, 29038, 28078, 28131, 28096, 28039, 28266, 28465, 28941, 28449, 28195, 25860, 24513, 25143, 23726, 21721, 19309, 17543, 16966, 17103, 16899, 17191, 16643, 17678, 15754, 19571, 7755, 477, 6841, 7106, 6250, 2329, 3998, 4704, 4508, 5191, 3305, 1420, 1323, 0, 215, 0, 54, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 594, 0, 2120, 0, 13833, 13681, 0, 4649, 1905, 4205, 3449, 4043, 3978, 4044, 3972, 3913, 4015, 3716, 3680, 1486, 4150, 0, 14486, 31819, 25768, 28316, 26900, 27610, 27338, 27321, 27595, 26588, 25716, 25761, 25067, 25451, 26122, 26641, 26861, 27089, 27423, 27414, 27437, 27596, 27648, 28257, 28333, 28463, 28403, 29344, 29690, 29107, 28810, 29037, 28849, 28226, 28367, 28652, 28070, 29660, 30388, 26944, 26018, 26410, 24836, 21708, 16641, 12826, 8740, 6170, 6965, 6483, 6908, 6374, 7290, 4583, 2585, 2477, 2089, 3312, 3431, 2872, 507, 0, 26, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 37, 0, 128, 0, 1528, 5901, 7786, 7316, 8174, 6533, 13726, 25104, 26446, 25638, 26406, 27600, 29877, 28008, 35579, 16060, 0, 2657, 377, 912, 2278, 0, 15009, 33388, 27637, 30232, 28364, 29350, 28856, 28880, 28854, 28843, 28844, 28854, 28828, 28884, 28705, 28593, 28764, 28798, 28885, 28889, 28806, 28806, 28717, 28783, 28674, 28804, 28933, 28694, 28702, 28312, 27998, 27960, 27563, 27259, 27790, 26905, 27280, 25377, 25822, 10013, 0, 1176, 0, 336, 0, 82, 0, 66, 0, 232, 0, 1863, 4253, 3454, 3985, 3463, 4182, 2904, 6755, 9203, 7581, 8596, 8042, 2946, 0, 332, 0, 91, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 242, 0, 858, 0, 7428, 18935, 18860, 18928, 25402, 28492, 35530, 16766, 0, 3957, 2268, 2396, 4676, 0, 16819, 36721, 30534, 33797, 31748, 33419, 30374, 28115, 28892, 28349, 28433, 28356, 28539, 28460, 28554, 28498, 28676, 28720, 28789, 28770, 28919, 29035, 28959, 29080, 29082, 28882, 29052, 28859, 29239, 28740, 29585, 23774, 11079, 8811, 3615, 0, 443, 0, 127, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 38, 0, 596, 2862, 3569, 4378, 5144, 5204, 5547, 5845, 2859, 487, 510, 0, 184, 0, 446, 0, 1427, 0, 12578, 33110, 25484, 29240, 32131, 27171, 25208, 25750, 25971, 29455, 14299, 0, 14681, 28909, 25106, 27016, 25878, 26639, 25980, 27306, 28443, 27859, 27958, 27646, 27392, 26931, 26545, 26361, 26081, 26097, 25936, 25902, 25994, 25604, 25973, 27028, 28262, 28588, 28486, 28727, 28534, 28639, 28395, 28449, 28849, 28796, 29450, 29431, 30470, 31587, 31037, 29557, 28653, 29092, 28110, 27939, 28226, 27968, 28275, 27761, 28671, 27025, 30350, 18575, 883, 360, 0, 126, 0, 8, 0, 0, 0, 1, 0, 9, 0, 35, 0, 255, 438, 301, 405, 357, 651, 287, 0, 35, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 35, 0, 310, 664, 4701, 15695, 25697, 25097, 33753, 16064, 0, 5800, 3238, 4916, 4151, 4604, 4502, 4558, 4627, 4754, 4810, 4487, 4101, 4064, 3824, 3674, 3724, 3683, 3734, 3656, 3758, 3417, 2552, 3360, 1744, 3990, 0, 14621, 33679, 28495, 29029, 28226, 28397, 28187, 28183, 28058, 27964, 28360, 27461, 29968, 25904, 35197, 16137, 0, 0, 13592, 33184, 26652, 29648, 27899, 27628, 28767, 26800, 31598, 13596, 0, 1668, 0, 466, 0, 28, 92, 0, 489, 0, 3828, 8447, 8232, 6621, 2565, 1078, 0, 363, 154, 0, 16, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 334, 0, 3043, 9046, 10904, 11362, 11369, 11075, 10522, 11023, 11238, 12980, 14080, 14337, 14221, 11361, 10370, 5262, 1273, 1187, 0, 202, 0, 48, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 40, 0, 135, 0, 1452, 5426, 6281, 6820, 6495, 6989, 3874, 1616, 1966, 4374, 3583, 11795, 21859, 22676, 26326, 26248, 27645, 28550, 29040, 29282, 29825, 30524, 30934, 31210, 30944, 31399, 30583, 32173, 27234, 23740, 26296, 25422, 25836, 17379, 15588, 16929, 18046, 18335, 22502, 10920, 0, 1253, 0, 356, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 124, 0, 433, 0, 3355, 6787, 4482, 4978, 3994, 3017, 3011, 3108, 3524, 2556, 4445, 627, 12802, 22599, 17737, 13988, 9708, 8479, 3644, 2876, 2089, 1021, 0, 126, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 157, 0, 547, 0, 4559, 11109, 9241, 10012, 10816, 14745, 14750, 17001, 21839, 23405, 25547, 26805, 23183, 20108, 17384, 9655, 7137, 8336, 8999, 9404, 9305, 9160, 8756, 8874, 7914, 5492, 4540, 3845, 2799, 4100, 1954, 0, 246, 0, 71, 0, 14, 0, 0, 0, 0, 0, 4, 0, 20, 0, 69, 0, 623, 1714, 1487, 1635, 2017, 2053, 2062, 1766, 2356, 1318, 0, 818, 3589, 7071, 9258, 11015, 11563, 12002, 12462, 13058, 14415, 15391, 16222, 16701, 16209, 17277, 12771, 7798, 7152, 5203, 5464, 5338, 6735, 6192, 4857, 5358, 5001, 5377, 4844, 5818, 2633, 0, 1844, 2829, 2763, 2966, 3145, 3042, 3298, 2609, 2004, 1375, 0, 3520, 14640, 21091, 17331, 7914, 4444, 1938, 135, 2201, 1832, 2756, 1190, 0, 65, 0, 6, 17, 0, 105, 0, 1021, 3239, 4086, 4380, 4840, 5293, 5170, 5198, 5243, 5106, 5413, 4357, 2749, 939, 0, 88, 0, 0, 230, 345, 789, 1855, 1922, 2100, 2101, 2924, 4213, 2555, 314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 232, 1813, 4228, 5072, 4808, 5066, 4696, 5312, 4138, 7957, 11701, 9716, 11454, 6017, 71, 184, 0, 66, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 52, 0, 188, 0, 1379, 2408, 1709, 1934, 2396, 3512, 3274, 2915, 3974, 4171, 4117, 2102, 0, 117, 0, 0, 440, 723, 2268, 4388, 4639, 4634, 3984, 1313, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 114, 0, 400, 0, 3278, 7799, 6982, 7941, 7847, 8725, 7721, 10850, 13581, 10742, 16475, 19671, 18221, 18858, 17800, 17377, 17592, 17616, 18744, 13171, 3615, 5519, 10141, 10675, 10292, 9694, 10115, 10573, 10441, 10512, 10464, 10503, 10507, 9661, 3423, 0, 949, 155, 28, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 51, 0, 235, 0, 1251, 467, 5487, 11977, 16407, 23321, 24567, 25379, 26023, 27241, 29481, 30340, 31314, 32582, 32075, 31723, 31235, 31451, 31249, 31528, 31060, 31973, 28890, 24602, 22450, 18579, 18230, 18450, 17682, 16721, 16504, 15009, 14405, 12995, 11334, 12249, 8707, 2686, 67, 29, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 36, 50, 1199, 1141, 2317, 3277, 3659, 4744, 4411, 4487, 4618, 4235, 5077, 2251, 0, 279, 0, 79, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 53, 0, 176, 0, 1489, 3578, 2147, 3157, 2676, 1540, 2159, 2861, 1143, 0, 0, 549, 0, 5292, 13149, 12478, 13024, 14064, 13246, 15033, 6674, 0, 828, 0, 220, 0, 0, 138, 144, 1014, 1773, 1530, 1445, 1017, 1077, 1261, 1301, 1311, 1277, 1344, 1219, 1469, 650, 0, 80, 0, 22, 0, 14, 0, 48, 0, 136, 0, 1730, 4515, 3202, 4617, 689, 5239, 15984, 14961, 16243, 21597, 25367, 26862, 27130, 26911, 26499, 25801, 23903, 20123, 18598, 18133, 18235, 19001, 19287, 17590, 16869, 15407, 13840, 14491, 13870, 14735, 13297, 16070, 7088, 0, 834, 0, 1440, 401, 0, 40, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 491, 663, 951, 2261, 2706, 4210, 5857, 6332, 5859, 5336, 5830, 5412, 5585, 5560, 5027, 4929, 4897, 4989, 4807, 5150, 4473, 6462, 6623, 3978, 3837, 4151, 3244, 3099, 3698, 4332, 4719, 1999, 284, 0, 10, 0, 0, 10, 0, 75, 99, 0, 100, 0, 314, 0, 2139, 2092, 0, 306, 0, 49, 28, 0, 582, 1310, 702, 1436, 2141, 2077, 2139, 2087, 2144, 2062, 2212, 1695, 923, 776, 208, 0, 18, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 18, 0, 62, 0, 697, 2686, 3483, 3738, 3773, 3916, 3724, 4063, 1641, 0, 192, 0, 55, 0, 11, 0, 0, 0, 0, 3, 0, 39, 0, 362, 1002, 2248, 1020, 5882, 9770, 7157, 5982, 4484, 4804, 4214, 3444, 3156, 2777, 2903, 3333, 2965, 2391, 1759, 1146, 266, 0, 22, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 34, 0, 134, 0, 1035, 2491, 4233, 3395, 2010, 4149, 7376, 11064, 14194, 15596, 16779, 18514, 18459, 18116, 20589, 20147, 19912, 19419, 19425, 21476, 21463, 21927, 19397, 18794, 17565, 16035, 14851, 14029, 14009, 13892, 13633, 14294, 12991, 15639, 6922, 0, 859, 0, 246, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 66, 0, 306, 0, 1393, 0, 8807, 17664, 15583, 18046, 17929, 18944, 19735, 19145, 21651, 24039, 23365, 23626, 23620, 23345, 24504, 25474, 24808, 25484, 23978, 21478, 19954, 21518, 19768, 20072, 24272, 21980, 25421, 14635, 3013, 6724, 2320, 0, 4300, 2645, 0, 335, 0, 103, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 200, 0, 699, 0, 5784, 13786, 11895, 12375, 12035, 11809, 13333, 16274, 17591, 18410, 19097, 19828, 19180, 20742, 21556, 22010, 23512, 24802, 26468, 26578, 27274, 27319, 28312, 29597, 30434, 29912, 28814, 29426, 30870, 31911, 30947, 31923, 29374, 31156, 15825, 505, 0, 10251, 21294, 17713, 19801, 18092, 20107, 16936, 24077, 12977, 0, 1409, 0, 891, 3157, 2830, 7670, 11990, 5299, 2790, 3402, 3788, 6532, 5969, 12185, 19997, 22061, 23564, 20789, 13864, 10339, 11727, 11149, 11029, 10229, 10019, 5024, 2878, 3033, 647, 262, 0, 39, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 71, 0, 222, 0, 3075, 5438, 3651, 5225, 1233, 5469, 14403, 12904, 19277, 26289, 27818, 27676, 29292, 24888, 18275, 18702, 18030, 18515, 17978, 18779, 17398, 20112, 11300, 2963, 5837, 4248, 4567, 4151, 1645, 0, 183, 0, 52, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 62, 0, 235, 0, 1644, 2835, 3581, 2939, 879, 1306, 1617, 500, 2833, 0, 13962, 30476, 24480, 26823, 18833, 16324, 12337, 6939, 7873, 7286, 3158, 0, 320, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 304, 0, 1063, 0, 8491, 18564, 14432, 18957, 21814, 20053, 15305, 15139, 15610, 18483, 19317, 25280, 31834, 30884, 32395, 30464, 27880, 24504, 13318, 7993, 9081, 8272, 8144, 7817, 7180, 4849, 1870, 0, 61, 0, 17, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 47, 0, 193, 0, 1390, 3077, 7626, 13357, 15781, 17070, 17057, 16266, 15762, 16624, 15430, 13131, 13547, 15334, 14542, 15407, 8053, 2322, 4180, 3885, 4604, 4956, 5243, 5330, 5221, 5385, 5881, 5857, 5744, 5487, 4802, 3653, 1035, 0, 101, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 20, 0, 97, 0, 322, 0, 2888, 7922, 6826, 9563, 10197, 9007, 10012, 9728, 10888, 11126, 11108, 9760, 9438, 7117, 6605, 4905, 10697, 16934, 16955, 20941, 22128, 24583, 27293, 29918, 30316, 30763, 30894, 30987, 30716, 31269, 30215, 32357, 25090, 15415, 12293, 9336, 9772, 8502, 8153, 7323, 5495, 4174, 3493, 3246, 2885, 2773, 1254, 0, 158, 0, 43, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 158, 477, 1835, 962, 5167, 10071, 9790, 10475, 10133, 10348, 10180, 10365, 10025, 11620, 15569, 12009, 7850, 8291, 8947, 9660, 10035, 10370, 10594, 10116, 9106, 8011, 6747, 6896, 6583, 6086, 5749, 4872, 5738, 2423, 0, 294, 0, 84, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 0, 370, 0, 1304, 0, 10915, 27192, 26155, 27785, 27515, 28944, 26540, 25427, 23119, 22610, 22659, 22991, 22004, 21243, 21987, 20817, 20475, 19753, 19761, 19555, 19298, 19225, 18757, 17821, 17634, 17476, 16628, 12636, 10868, 12694, 11325, 9619, 3188, 0, 349, 0, 101, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 130, 0, 450, 0, 3432, 6626, 4199, 6090, 5053, 1463, 0, 1085, 3127, 4107, 6660, 9248, 10110, 10665, 12122, 12112, 11790, 13148, 14061, 13581, 10033, 2729, 0, 259, 0, 73, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 104, 0, 346, 0, 3144, 8727, 6790, 8414, 9434, 8985, 6673, 5944, 3693, 6328, 13606, 17574, 20540, 21582, 19817, 16586, 11670, 7902, 8840, 8706, 8182, 9681, 4326, 0, 535, 0, 153, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 0, 92, 295, 322, 261, 577, 2804, 3816, 3801, 3398, 4336, 2331, 9263, 17683, 16775, 17817, 18013, 17019, 17538, 13146, 9150, 8924, 9811, 4513, 0, 567, 0, 156, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 149, 0, 531, 0, 4247, 10052, 10194, 7232, 716, 18, 0, 2, 85, 229, 0, 1441, 0, 5000, 0, 22866, 21195, 0, 11166, 9357, 11385, 9915, 7570, 6251, 5062, 3811, 4060, 1161, 0, 106, 0, 34, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 0, 158, 659, 518, 802, 0, 4002, 10840, 12173, 13472, 14129, 15230, 15290, 15951, 16604, 17162, 16242, 13773, 13419, 7399, 1044, 519, 0, 97, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 13, 0, 27, 502, 4908, 5733, 6682, 11241, 8609, 1983, 0, 1012, 1835, 4558, 6486, 7988, 9383, 9858, 9896, 9755, 9875, 9794, 9893, 9733, 10015, 9454, 11339, 13539, 12872, 11888, 10826, 10515, 9829, 9399, 8741, 8069, 8280, 6749, 1748, 0, 153, 0, 44, 0, 10, 0, 0, 0, 0, 0, 0, 27, 0, 131, 0, 457, 0, 3718, 8442, 7106, 11287, 14954, 15435, 14596, 14421, 14348, 14575, 14107, 14989, 13209, 19237, 26504, 25589, 26607, 26873, 26905, 25026, 20788, 16907, 11798, 10093, 4166, 0, 510, 0, 141, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 54, 0, 179, 0, 1518, 3443, 853, 0, 107, 980, 1152, 1152, 1104, 3504, 5863, 12850, 17958, 18624, 20353, 21910, 21201, 18547, 17094, 16906, 9082, 1240, 1146, 0, 210, 0, 45, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 135, 0, 495, 0, 3968, 9704, 11533, 14497, 15527, 20109, 13547, 1840, 3892, 10457, 12599, 14259, 14268, 12075, 11592, 11620, 10962, 10941, 10853, 10624, 10818, 10498, 11071, 10032, 12093, 5349, 0, 664, 0, 190, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 0, 0, 998, 8574, 12382, 11983, 7243, 3557, 7770, 6567, 3095, 1068, 2105, 3101, 6367, 6434, 6657, 10555, 11470, 12138, 11916, 11994, 12007, 11909, 12136, 11346, 10353, 10435, 9936, 10101, 10110, 10256, 8925, 7043, 2406, 0, 269, 0, 75, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0);


--  Datos de 1 a 16
--    type t_reg_datos is array (0 to 32783) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (20281, 19442, 16957, 15142, 15412, 15158, 15446, 15015, 15796, 13576, 13213, 14746, 14148, 13681, 14541, 16329, 16067, 17112, 17673, 17879, 17338, 16618, 17513, 17677, 18974, 19412, 19299, 20713, 20716, 21630, 19675, 17264, 17171, 15561, 14850, 14784, 14268, 13055, 12547, 12652, 15122, 16961, 15195, 15539, 15896, 16354, 18070, 17031, 15867, 16308, 15920, 16433, 15532, 18360, 21149, 20358, 20118, 20773, 18637, 15919, 16950, 15582, 14798, 14490, 13714, 12949, 12545, 12596, 14971, 15943, 14995, 15356, 15244, 15672, 15149, 16057, 12456, 12160, 14705, 14746, 17536, 19683, 20632, 19339, 18951, 18961, 18166, 16160, 14775, 13998, 13819, 14098, 13968, 14087, 13927, 14190, 13695, 15172, 15826, 15349, 15793, 15411, 15282, 15425, 13628, 10017, 13746, 17765, 18410, 19097, 18160, 18291, 18266, 18194, 16299, 14385, 14564, 14430, 14794, 15266, 14333, 13756, 13479, 13309, 14106, 14906, 15300, 15144, 15461, 16010, 15456, 16309, 13637, 10992, 11725, 11282, 11449, 11483, 11226, 11807, 10600, 14305, 16406, 15236, 13275, 13058, 15040, 13489, 14385, 13898, 13520, 14624, 14786, 15443, 16125, 15897, 16159, 16090, 16773, 16294, 17475, 13735, 13670, 18340, 18214, 19152, 18688, 18990, 19240, 18986, 18450, 16352, 15067, 14897, 14771, 13998, 13388, 13457, 13339, 13298, 13285, 13327, 13245, 13388, 13092, 14315, 16772, 14728, 11917, 10636, 15085, 21140, 22611, 22406, 19945, 18489, 18989, 17788, 16992, 14503, 12555, 13098, 12361, 12425, 12993, 13356, 13007, 12966, 16652, 20103, 14402, 12960, 15909, 16334, 17999, 14797, 12790, 12737, 15005, 21705, 24848, 24482, 20347, 18059, 18770, 18263, 18819, 18002, 19501, 14603, 9666, 13565, 13866, 12085, 13051, 17623, 19252, 14209, 14067, 15731, 15216, 18963, 15817, 11225, 14981, 17980, 20281, 24541, 22807, 20467, 19093, 17833, 17734, 17626, 14109, 11981, 12690, 12902, 14158, 12030, 12482, 11230, 12450, 15248, 18058, 13732, 10762, 13912, 12626, 13377, 12833, 13384, 12527, 15303, 19022, 17438, 14309, 12046, 12024, 11579, 10825, 10179, 9118, 8125, 2635, 0, 255, 65, 1114, 3226, 7181, 4937, 4904, 5229, 2274, 2739, 3468, 3943, 3801, 7301, 6678, 7174, 10900, 8869, 8498, 8904, 9335, 9643, 7035, 3477, 966, 593, 639, 616, 637, 614, 646, 432, 0, 920, 1607, 2215, 1551, 3975, 8143, 8214, 10267, 9741, 7938, 10131, 10187, 7457, 5714, 6561, 8137, 8270, 7601, 2265, 0, 225, 0, 67, 0, 14, 0, 26, 0, 137, 0, 490, 0, 3741, 7569, 6772, 8447, 7694, 8055, 7896, 7942, 7960, 7852, 8708, 10921, 4059, 0, 455, 0, 149, 0, 108, 0, 273, 0, 1795, 1923, 0, 581, 0, 2464, 5584, 6427, 7625, 6219, 6980, 7178, 7515, 9055, 9759, 8363, 8337, 3322, 0, 396, 0, 113, 0, 22, 0, 0, 5, 0, 25, 0, 85, 0, 1129, 5119, 7333, 7720, 7425, 6328, 7226, 7642, 8519, 10360, 9287, 10455, 4203, 0, 502, 0, 146, 0, 29, 0, 0, 0, 0, 22, 0, 107, 0, 365, 0, 3117, 7916, 6425, 6725, 6224, 6632, 7095, 7462, 9068, 9327, 9414, 9186, 9628, 8807, 10461, 4833, 0, 1652, 748, 0, 56, 0, 0, 79, 0, 1299, 5605, 7450, 7420, 8089, 7137, 7347, 7928, 7175, 8053, 8066, 7902, 6757, 1869, 0, 216, 0, 165, 0, 1621, 6307, 2332, 684, 2183, 0, 958, 48, 3849, 7098, 6110, 6637, 6305, 6562, 6266, 7096, 8173, 7923, 8830, 8909, 8653, 7891, 6772, 2250, 0, 0, 1635, 7379, 8126, 8533, 10605, 7486, 1583, 3259, 5942, 7265, 9388, 10075, 10243, 10946, 13124, 15126, 11046, 7483, 9598, 10056, 10725, 9051, 7840, 7345, 7244, 6372, 3654, 2900, 3028, 2991, 2975, 3060, 2833, 3762, 6458, 10692, 11310, 10331, 10642, 12155, 15508, 15761, 16054, 13437, 11339, 14072, 13996, 13475, 12873, 11615, 12032, 12772, 10522, 7813, 8735, 8864, 8034, 11356, 15652, 11520, 7766, 9196, 10968, 13339, 11543, 9800, 11402, 15953, 17335, 17562, 17249, 15480, 16118, 15775, 15985, 15834, 16004, 15238, 12837, 13847, 12237, 10779, 9816, 11283, 14596, 15024, 13224, 8358, 11357, 13157, 13102, 14028, 11838, 15129, 18273, 18704, 20247, 19379, 17872, 16548, 16950, 16816, 14881, 15317, 15546, 15735, 14612, 14881, 14038, 11290, 11287, 13466, 14409, 16901, 14288, 10132, 11380, 10918, 10863, 11461, 9962, 15185, 20963, 20440, 20258, 19894, 19252, 16721, 17812, 14863, 14061, 16449, 16516, 15066, 13806, 13506, 10511, 11441, 14931, 16351, 18347, 16891, 14023, 17214, 17828, 17517, 14797, 11401, 17224, 20947, 20630, 21565, 21323, 20805, 20329, 19229, 16600, 14057, 14093, 14225, 14196, 14227, 14176, 14268, 14082, 14738, 16248, 17976, 16379, 13947, 16160, 16820, 17745, 15421, 9689, 14072, 19190, 19611, 20900, 20795, 20884, 20767, 19269, 18155, 15030, 13536, 14480, 14349, 14608, 14567, 15113, 14789, 13605, 15000, 18023, 18708, 18917, 16311, 16784, 19585, 18798, 20182, 16139, 12803, 13937, 13105, 14026, 12562, 17046, 21469, 18214, 15494, 14608, 14335, 15595, 15708, 14321, 15321, 15338, 14314, 14613, 17024, 18941, 18795, 16204, 16422, 19190, 18850, 20022, 15168, 11334, 17152, 19513, 19939, 21029, 20792, 20773, 20717, 17569, 16641, 16440, 16247, 16519, 16473, 15031, 14039, 14823, 14592, 14811, 14553, 14947, 14206, 16551, 18821, 19041, 18723, 14112, 11088, 15502, 19163, 18715, 19994, 20587, 20987, 19883, 17590, 16950, 15847, 14356, 15459, 16560, 15901, 15070, 13276, 11730, 13861, 15860, 17149, 18856, 18175, 17988, 18517, 18748, 19746, 14428, 10815, 16516, 19356, 19377, 19850, 19812, 19905, 19801, 19949, 19712, 20165, 18572, 16401, 17048, 14936, 15206, 15173, 14653, 16057, 17998, 18218, 15804, 16545, 18333, 18704, 19847, 15051, 9722, 16100, 19637, 19678, 20378, 19918, 20081, 19661, 18705, 16859, 15487, 14896, 14466, 14827, 15808, 15330, 17227, 14345, 13736, 17507, 17594, 18899, 18851, 18930, 18910, 18884, 18956, 18811, 19247, 19599, 20003, 20339, 20718, 20920, 20182, 19225, 17674, 17306, 17460, 17100, 16879, 16271, 16435, 16475, 16062, 16113, 17085, 18384, 20138, 21258, 20815, 20745, 19765, 21504, 18647, 15977, 18963, 20229, 21507, 22091, 22165, 21312, 20594, 20249, 20086, 18347, 17225, 17521, 17407, 17412, 17514, 17241, 18278, 19862, 20198, 21729, 23169, 23408, 22883, 21507, 22092, 22299, 21487, 20842, 20550, 21584, 21844, 21899, 21064, 20738, 20364, 18778, 17499, 17717, 17025, 16836, 16756, 16831, 17719, 16325, 15754, 16647, 16994, 18597, 19550, 18348, 18831, 18222, 20358, 15940, 11093, 12523, 11935, 12015, 12410, 11312, 15033, 17790, 16113, 16788, 13767, 13143, 15471, 15399, 15222, 14088, 12380, 10638, 13166, 15917, 16319, 17270, 16409, 16357, 15903, 18089, 13695, 11388, 11669, 13521, 17531, 18329, 17603, 16121, 17036, 15898, 16002, 13961, 12099, 13014, 14431, 14699, 15430, 13642, 11681, 12209, 12095, 11880, 12510, 11113, 15743, 20361, 20093, 19120, 17094, 20220, 20611, 19873, 20153, 20818, 20987, 20723, 20660, 18043, 16835, 16638, 17312, 18536, 18256, 18722, 18593, 18417, 18077, 19014, 20006, 20503, 21940, 21918, 21666, 21331, 21651, 21623, 20151, 20580, 20505, 19919, 19328, 19539, 20230, 19988, 20130, 20013, 20156, 19934, 20203, 17684, 16194, 16945, 17566, 16462, 16662, 18657, 19169, 20838, 20501, 20893, 20445, 20656, 20855, 19221, 19501, 19071, 18286, 17645, 18226, 19728, 19857, 20516, 19829, 17174, 15080, 15992, 16471, 15062, 14414, 13557, 13869, 14218, 15119, 17115, 18691, 18914, 18580, 18709, 18616, 18724, 18551, 18863, 18133, 18364, 15830, 13589, 15120, 14713, 15246, 16053, 15521, 15152, 15590, 15633, 15438, 15363, 14548, 13330, 13065, 14661, 15036, 17719, 18408, 18015, 20394, 20470, 21159, 20305, 19571, 19192, 19492, 19246, 16803, 17856, 18577, 18772, 18754, 18662, 19031, 18623, 19072, 18914, 18941, 19025, 18804, 19273, 17786, 16972, 18806, 19569, 20623, 20650, 19968, 19779, 18803, 18441, 17596, 18267, 19323, 17268, 17503, 18558, 18968, 20062, 19570, 19947, 19936, 20530, 20483, 18232, 17304, 16281, 16731, 17839, 19169, 17754, 18701, 19890, 21362, 20445, 19595, 20930, 19705, 20613, 20545, 20641, 20571, 20645, 20532, 20743, 20109, 20049, 21585, 21041, 21547, 20597, 19792, 19844, 18925, 18633, 19976, 20369, 18756, 19835, 20773, 22396, 21882, 21399, 22636, 21728, 21979, 22119, 21897, 22238, 21543, 20891, 20668, 20976, 21683, 21640, 21151, 22192, 21458, 19742, 20137, 19120, 18131, 18930, 19300, 19174, 19329, 19066, 19537, 18628, 21372, 22940, 22010, 23210, 22055, 23772, 24015, 22753, 22965, 22504, 22424, 22446, 22208, 22751, 22751, 22768, 21805, 21795, 21022, 19172, 20004, 20124, 21045, 22316, 21595, 20749, 20764, 22691, 23159, 21718, 21988, 23110, 22205, 23220, 24502, 23425, 24121, 23879, 23631, 23717, 23640, 23736, 23589, 23865, 22931, 21683, 21929, 22501, 21997, 21229, 22531, 23140, 22670, 22846, 22199, 22367, 21840, 21632, 22843, 23079, 22151, 22119, 23459, 23930, 24182, 22964, 22752, 22965, 22415, 23357, 23692, 22440, 22035, 21641, 21550, 22266, 22083, 22797, 23654, 23153, 22047, 22150, 22662, 22496, 22577, 22540, 22546, 22567, 22583, 23494, 24453, 24971, 23851, 23081, 23220, 22914, 22993, 22507, 22303, 22661, 22018, 21586, 22611, 21584, 23130, 24542, 22856, 22155, 22283, 22374, 23379, 22852, 22123, 23380, 22802, 23146, 23936, 24669, 25235, 24608, 24078, 23536, 22986, 22137, 21445, 22548, 23201, 23025, 23122, 23049, 23124, 23024, 23173, 22101, 20162, 20176, 21106, 21454, 21176, 21326, 21634, 21672, 22184, 22296, 23203, 23916, 23891, 22567, 21314, 20336, 20060, 20993, 21167, 21249, 21164, 21288, 20632, 20546, 20042, 21467, 23147, 21406, 19880, 19827, 20252, 21058, 20462, 19998, 21131, 20520, 19988, 20137, 20057, 20108, 20072, 20112, 19919, 19052, 18484, 18284, 18523, 18777, 17661, 17295, 16575, 17365, 18433, 20520, 20103, 17864, 18706, 19168, 20000, 20184, 19944, 19534, 18360, 19710, 21108, 21214, 22027, 21600, 21043, 19431, 18358, 17862, 17880, 17746, 17216, 17310, 16892, 16206, 16297, 16576, 16563, 16549, 16614, 16468, 16755, 16172, 17987, 19090, 18354, 18165, 19711, 19827, 18805, 20217, 19896, 18950, 18080, 17749, 17409, 17081, 16151, 15824, 14641, 14602, 15526, 15361, 14517, 15111, 14635, 16489, 17884, 16678, 17309, 17983, 19085, 18465, 18285, 17317, 18171, 18945, 18097, 19197, 19909, 19158, 18823, 18776, 19008, 18520, 19528, 16160, 12615, 13650, 13447, 14573, 14711, 14870, 16331, 16913, 16365, 16170, 17020, 18034, 17324, 16363, 15948, 17105, 18052, 18041, 18207, 18521, 17600, 16925, 16203, 15367, 15007, 14359, 14672, 14163, 13598, 13649, 13702, 14018, 14805, 14622, 14979, 15816, 15701, 16476, 17066, 16907, 16963, 16981, 16876, 17154, 17083, 18845, 19087, 17665, 18386, 16635, 15991, 14861, 14353, 15129, 14246, 14322, 13996, 14161, 14402, 14842, 14656, 14770, 15819, 15910, 16360, 15903, 16336, 15398, 11657, 14541, 18052, 17135, 17478, 17790, 18248, 17843, 17523, 16147, 15325, 13228, 11507, 13367, 13622, 13703, 13553, 13815, 13306, 14774, 14717, 12966, 13157, 14140, 15909, 16019, 16663, 13971, 15076, 18813, 18232, 19076, 18629, 17955, 17800, 17424, 17025, 15942, 15830, 15862, 15995, 15034, 14499, 14539, 14189, 14973, 15755, 14871, 12697, 12235, 12300, 13476, 15618, 15720, 16529, 14521, 15926, 18815, 17862, 18357, 18067, 18263, 18083, 18275, 17001, 15817, 14654, 13660, 14348, 13337, 14686, 12378, 12461, 15777, 15419, 13850, 13204, 14400, 14703, 16901, 17308, 14988, 12878, 16271, 18966, 18395, 19010, 18285, 17857, 17803, 17834, 18601, 17024, 15687, 16041, 16588, 16871, 15002, 14425, 14693, 15134, 15743, 15512, 15672, 15517, 15720, 15354, 16740, 18778, 15919, 16679, 19339, 18116, 17912, 18139, 17935, 17791, 17812, 18008, 16714, 15010, 16251, 16784, 16585, 15701, 15116, 14448, 15071, 16740, 17171, 17107, 16663, 17124, 17614, 18261, 18404, 18764, 18443, 18376, 19021, 17875, 17218, 17698, 17424, 17199, 17121, 17164, 17100, 17214, 17007, 17419, 16079, 14938, 16210, 16952, 17556, 16829, 15975, 16347, 17029, 17410, 17629, 18323, 18434, 18004, 18807, 18448, 17900, 18317, 18301, 18236, 17581, 18060, 17616, 16960, 17066, 17034, 16113, 15246, 15743, 16570, 15383, 15784, 17132, 16029, 16049, 16903, 17405, 17475, 17765, 17661, 17717, 17680, 17716, 17660, 17860, 18320, 18572, 18097, 18032, 17589, 15921, 14980, 15054, 15033, 15140, 16526, 13353, 10618, 15439, 16819, 16681, 16398, 15656, 16736, 16983, 17792, 19086, 17095, 16842, 18838, 17748, 17796, 17886, 18139, 18496, 18178, 18269, 17407, 16940, 17342, 17239, 15912, 14954, 15222, 15109, 15136, 15184, 15029, 15598, 16415, 17089, 17636, 18048, 18791, 17820, 17721, 18177, 17058, 16788, 17769, 18406, 18055, 17898, 16939, 16416, 15497, 13603, 14502, 14278, 15185, 14619, 13733, 15205, 15537, 16479, 15931, 15313, 16704, 17438, 17835, 17097, 15877, 14594, 16431, 18264, 17037, 17322, 17181, 17167, 17351, 16930, 17808, 15045, 12894, 12793, 13546, 14110, 12176, 10790, 13836, 17425, 15847, 15136, 13414, 13862, 14867, 15067, 16260, 16048, 14548, 16361, 18112, 17303, 17213, 17507, 17628, 17411, 17414, 16276, 16212, 15062, 13954, 12458, 12290, 12812, 10822, 13126, 16335, 17302, 15525, 14296, 14607, 14526, 14441, 14723, 14086, 16224, 18269, 17334, 17375, 17076, 17724, 17604, 17275, 17266, 17348, 15843, 13985, 15081, 14478, 14844, 13655, 13911, 16738, 16893, 17977, 16885, 15335, 16273, 16740, 17285, 18492, 18491, 18002, 18105, 18475, 18117, 17811, 17633, 17935, 17581, 17696, 16669, 16406, 17296, 16970, 17139, 17051, 17086, 17081, 17209, 18090, 16558, 14379, 13579, 15512, 17210, 17202, 14957, 15364, 18369, 18080, 18562, 18350, 18228, 18611, 18019, 17835, 17374, 16867, 16650, 15941, 16107, 16678, 16272, 16083, 15410, 16690, 17332, 16519, 15884, 15363, 15054, 16548, 17279, 16660, 15713, 16437, 18564, 17841, 18216, 17994, 18153, 17990, 18223, 17192, 16175, 16085, 16095, 16032, 16423, 16627, 16036, 15876, 16265, 16877, 16682, 16139, 16147, 16167, 17701, 18223, 17249, 18594, 19373, 19811, 19952, 19605, 19665, 18873, 18260, 17844, 18564, 17596, 16249, 16597, 16242, 16554, 16483, 15998, 15924, 15965, 15802, 15844, 15857, 15783, 15947, 15608, 16681, 17591, 17964, 19396, 19880, 19763, 19132, 19458, 19256, 17883, 17782, 18291, 17106, 15893, 17079, 17446, 17765, 17078, 16026, 15909, 16355, 17300, 17428, 16956, 17340, 18382, 18010, 18212, 18405, 18846, 19310, 19805, 19449, 19257, 18809, 18539, 18562, 17917, 17967, 17933, 17914, 17995, 17824, 18173, 17054, 15949, 15693, 15648, 16941, 17157, 16957, 17892, 18463, 18091, 18349, 18712, 18970, 18792, 18313, 18964, 19168, 19168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 75, 0, 327, 0, 2770, 6270, 5629, 0, 10661, 24447, 17811, 19006, 19355, 19646, 19980, 20235, 20679, 21353, 21611, 21753, 21756, 21986, 22034, 22426, 22159, 21898, 22147, 21543, 22148, 22492, 24410, 26015, 25737, 25488, 26324, 24583, 28178, 16344, 4833, 8428, 6593, 6552, 7611, 8549, 4108, 632, 3266, 2319, 0, 324, 0, 91, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 166, 0, 576, 0, 8443, 8730, 7098, 22821, 26982, 26424, 26509, 26703, 26127, 27444, 22951, 18922, 21343, 20781, 21230, 21519, 22905, 23671, 23448, 23399, 23198, 22542, 22695, 22738, 25128, 27074, 25322, 25960, 23176, 24912, 12790, 3700, 8316, 7956, 8945, 4867, 5206, 5986, 5111, 3746, 3574, 1577, 0, 196, 0, 54, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 174, 0, 554, 0, 5199, 12994, 1916, 5313, 22010, 27454, 27960, 27468, 27463, 26800, 23059, 21250, 21225, 20984, 19712, 19163, 19173, 18763, 18107, 17169, 17859, 18692, 20813, 21527, 24366, 26665, 25340, 28365, 30588, 30068, 30126, 30475, 29568, 31511, 25536, 21279, 16147, 7399, 4923, 311, 75, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 294, 0, 1040, 0, 8931, 21965, 16425, 12226, 21437, 30903, 29576, 30227, 29736, 28170, 26731, 27242, 26845, 27329, 26553, 28018, 23431, 19770, 21580, 21012, 21954, 21957, 22336, 22771, 24640, 27616, 28873, 26922, 28504, 28949, 29880, 23396, 14565, 7326, 2179, 3496, 1657, 1788, 1404, 1757, 811, 0, 236, 266, 120, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 35, 0, 93, 765, 9327, 12286, 13119, 24147, 29733, 30656, 31220, 30030, 32372, 27234, 37030, 10691, 13284, 36475, 33755, 17856, 0, 4576, 122, 1833, 1801, 1645, 1730, 3958, 2798, 2471, 2253, 5341, 0, 18031, 31694, 23601, 25727, 22468, 23920, 23467, 23181, 24253, 22038, 26537, 11743, 0, 1458, 0, 417, 0, 84, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 216, 0, 778, 0, 5941, 12045, 11512, 15774, 18464, 26572, 30758, 31092, 31141, 31175, 30307, 29069, 26263, 24898, 24061, 22585, 22786, 22689, 22605, 22975, 22125, 23882, 22341, 33055, 17070, 0, 4778, 1280, 4412, 1885, 5695, 0, 16400, 34338, 21858, 22097, 19843, 21733, 9119, 0, 1501, 0, 328, 0, 3008, 5137, 5295, 5962, 6283, 6140, 6914, 2769, 0, 322, 0, 59, 268, 2222, 3583, 3399, 3354, 3273, 3442, 3125, 3762, 1666, 0, 206, 0, 59, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 0, 353, 0, 1275, 0, 9351, 17532, 18463, 30582, 30982, 31375, 27701, 24183, 20862, 19427, 20510, 19734, 19898, 20062, 21080, 21131, 22754, 25385, 26120, 26485, 26731, 28236, 27219, 29519, 28584, 36394, 15409, 201, 545, 17031, 32934, 26218, 30123, 23444, 23860, 21479, 18098, 6727, 657, 2318, 1469, 1997, 1594, 2053, 876, 0, 111, 0, 31, 0, 1, 5, 0, 41, 0, 144, 0, 1311, 4248, 4409, 4212, 2587, 8190, 4959, 0, 678, 0, 194, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 173, 0, 558, 0, 4903, 13632, 10760, 12193, 4752, 14757, 26826, 24124, 22492, 17886, 20167, 19542, 19687, 19751, 19643, 19596, 19744, 19678, 19460, 19679, 21084, 21918, 21980, 22161, 22032, 22210, 21909, 22467, 21345, 24946, 28216, 29992, 30717, 32290, 24487, 20713, 13511, 2448, 2781, 6145, 10501, 8753, 5454, 2112, 4543, 5401, 5458, 5418, 4968, 5741, 2480, 0, 305, 0, 83, 0, 0, 34, 0, 152, 0, 1194, 2653, 2411, 1643, 111, 23, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 0, 336, 0, 1172, 0, 9465, 21532, 17930, 20160, 19409, 20137, 19972, 20464, 21598, 22190, 22062, 22117, 22121, 20881, 21115, 22280, 21191, 24536, 27609, 25388, 26336, 24396, 26775, 11514, 0, 5821, 5471, 7860, 4281, 4915, 6558, 5395, 5509, 5299, 6497, 1318, 2152, 5535, 3738, 4605, 4057, 4504, 3985, 4852, 2140, 0, 266, 0, 76, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 56, 0, 301, 0, 1097, 0, 7512, 10349, 7680, 17157, 20731, 20823, 17866, 19375, 18926, 18983, 18990, 18337, 17932, 18150, 18433, 20121, 22128, 20898, 21649, 21947, 20112, 20713, 19240, 22693, 25420, 24179, 24780, 24368, 24768, 24213, 25221, 22422, 20291, 12323, 10417, 16117, 16797, 6793, 0, 808, 0, 222, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 55, 0, 266, 0, 901, 0, 7292, 16404, 10411, 9532, 3061, 0, 333, 0, 100, 0, 1, 12, 0, 579, 3188, 3345, 3013, 4316, 6446, 9381, 2366, 2476, 10166, 6420, 1123, 46, 1847, 3623, 4741, 4817, 4994, 3087, 1195, 1408, 399, 0, 34, 0, 11, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 139, 0, 578, 0, 4213, 6953, 7073, 0, 10925, 29291, 27497, 30505, 29671, 29981, 29018, 29269, 28813, 29797, 27399, 35940, 16655, 0, 3612, 938, 3863, 2983, 4082, 3826, 3819, 3908, 3381, 4735, 4832, 3975, 4826, 5298, 4278, 3793, 3937, 3715, 4123, 3374, 4773, 1939, 11412, 21981, 21526, 21747, 24236, 11863, 343, 3829, 2984, 5373, 4990, 5905, 2233, 0, 213, 0, 0, 283, 0, 2525, 5830, 5616, 11457, 5155, 0, 632, 0, 190, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 142, 0, 1656, 951, 10110, 19968, 18014, 15332, 23704, 31568, 27623, 26932, 21899, 18646, 19994, 20518, 21417, 21528, 21757, 21255, 22268, 20146, 27157, 33304, 30704, 26523, 33761, 16065, 0, 6029, 3735, 6255, 3701, 6974, 0, 16898, 32178, 22989, 24782, 21653, 21318, 18871, 17965, 14925, 8906, 6678, 6643, 4879, 1576, 0, 165, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 220, 0, 745, 0, 6599, 18317, 17606, 17449, 11782, 9501, 14771, 18037, 19353, 19555, 21088, 22368, 22564, 22925, 22693, 24015, 25719, 26164, 26197, 26496, 26675, 25367, 23683, 23390, 22487, 24233, 24640, 26125, 25856, 31745, 14293, 0, 6574, 5039, 5609, 5498, 5927, 5360, 4792, 5041, 4818, 5118, 4621, 5580, 2466, 0, 306, 0, 87, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 201, 0, 739, 0, 6289, 7752, 10043, 25571, 29380, 27964, 25182, 23136, 22001, 22963, 23318, 25077, 28278, 30227, 28998, 28219, 29508, 30867, 31478, 31423, 31230, 31723, 30743, 32735, 26568, 23168, 26307, 25041, 26694, 32204, 23471, 8070, 6915, 7042, 6264, 4719, 2746, 1283, 1628, 1246, 387, 0, 38, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 303, 0, 1058, 0, 8665, 20427, 18094, 20105, 19299, 19518, 19531, 20414, 20859, 23993, 24168, 22039, 22384, 22058, 22078, 21939, 22915, 23723, 24363, 23347, 25561, 23895, 25455, 10384, 0, 1804, 11496, 25290, 21153, 24882, 12387, 4633, 5088, 548, 2366, 454, 0, 23, 0, 19, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 71, 0, 127, 0, 3120, 14620, 3123, 8736, 27861, 26540, 26940, 20617, 19423, 20666, 20358, 20788, 20514, 20586, 20632, 21010, 21447, 21598, 21847, 21762, 21614, 21712, 21684, 21135, 20056, 19449, 19770, 19304, 20149, 18562, 21759, 11908, 4748, 4570, 15122, 15759, 4210, 6259, 3188, 4389, 2948, 1357, 54, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 34, 0, 120, 0, 791, 791, 0, 120, 0, 34, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 156, 0, 441, 0, 4605, 13047, 416, 9381, 23311, 19751, 21691, 20611, 21200, 20879, 21086, 20781, 20851, 21069, 21268, 21521, 21502, 21463, 21414, 20808, 19842, 19758, 19531, 19245, 19774, 20196, 22417, 26060, 9373, 0, 2470, 4564, 5722, 6112, 6245, 3193, 2828, 3567, 2308, 1844, 2317, 438, 0, 17, 0, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 140, 0, 542, 0, 4467, 10177, 9820, 5704, 16159, 26542, 22104, 21286, 19370, 20456, 20122, 20834, 20865, 21868, 22682, 22687, 22418, 21763, 21901, 21942, 21823, 21634, 20678, 19560, 19803, 19547, 20109, 20072, 24002, 25830, 26170, 29641, 29740, 30008, 29619, 30295, 29047, 31468, 24898, 24278, 17019, 5217, 9596, 6269, 1721, 0, 144, 0, 27, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 208, 0, 726, 0, 5144, 7295, 0, 428, 0, 449, 0, 1211, 0, 9764, 22779, 19920, 21993, 21525, 22500, 22355, 22727, 22712, 22649, 22462, 22175, 22245, 23415, 24310, 23310, 25596, 26765, 26232, 25788, 23704, 16963, 7635, 6302, 7609, 7176, 6710, 6406, 7174, 5756, 7187, 2159, 2006, 3172, 0, 534, 0, 141, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 67, 0, 367, 0, 2527, 4719, 13051, 4192, 10784, 29093, 24098, 26087, 20160, 17323, 17202, 16831, 18728, 18935, 19739, 20509, 20471, 21245, 20590, 21306, 21444, 21458, 22101, 22409, 23052, 23038, 24725, 25449, 25467, 25105, 25918, 24354, 27546, 16493, 2581, 6881, 5338, 4850, 6118, 4775, 3875, 3289, 3763, 1595, 0, 195, 0, 55, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 177, 0, 626, 0, 5133, 11085, 6938, 10189, 20974, 26192, 24857, 25469, 25169, 25283, 25329, 24758, 22907, 21717, 21796, 21622, 20769, 19538, 18524, 17945, 17132, 18053, 17520, 21334, 23863, 25448, 23968, 28939, 16337, 0, 17037, 29176, 18510, 20774, 21296, 20770, 17421, 8941, 3959, 2282, 166, 27, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 86, 0, 295, 0, 3131, 3702, 137, 346, 0, 79, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 285, 0, 1000, 0, 8638, 21538, 16159, 13261, 21636, 29575, 27952, 27925, 26789, 25580, 23915, 23225, 23805, 24172, 23845, 24263, 24481, 22682, 21847, 22376, 21432, 21471, 22574, 22382, 23591, 23228, 26782, 29437, 27664, 27730, 28779, 30304, 30046, 30513, 29690, 31192, 28428, 33954, 15838, 0, 3759, 3016, 1805, 539, 1535, 0, 247, 0, 65, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 253, 0, 945, 0, 6519, 10420, 13944, 25681, 28057, 32194, 31111, 30982, 31465, 30255, 29709, 29825, 30064, 29389, 30761, 28172, 33372, 16262, 0, 4464, 2037, 3327, 1018, 283, 1589, 3123, 2313, 5910, 0, 15922, 28910, 21228, 24678, 21842, 20743, 17218, 15885, 5692, 0, 1890, 283, 9, 0, 0, 3, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 233, 0, 832, 0, 8584, 15103, 13898, 16241, 15719, 26192, 30702, 30147, 30385, 29296, 28610, 24131, 21064, 22914, 23700, 24064, 24287, 25235, 25568, 26515, 27110, 26742, 22008, 30960, 14769, 0, 4459, 2351, 3381, 3214, 2311, 5740, 0, 16484, 33165, 20601, 21438, 19858, 20597, 19805, 20928, 18981, 22838, 10127, 0, 1327, 0, 609, 0, 2378, 5308, 4453, 1633, 0, 191, 0, 43, 0, 0, 46, 0, 431, 916, 205, 0, 11, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 109, 0, 285, 0, 6813, 14298, 2704, 6514, 16818, 24501, 28628, 25815, 22844, 18460, 20331, 19622, 20177, 20028, 20077, 19546, 20887, 22736, 22753, 22866, 22753, 22907, 22645, 23405, 24383, 26457, 29972, 21105, 5804, 0, 8703, 20494, 17892, 24042, 25245, 19309, 21316, 9423, 73, 2624, 1142, 1863, 1111, 1456, 668, 2039, 1424, 0, 203, 0, 57, 0, 8, 0, 0, 12, 0, 40, 0, 529, 2310, 2902, 2807, 2791, 2903, 2651, 3183, 1411, 0, 175, 0, 50, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 444, 0, 1528, 0, 12570, 29134, 21075, 21415, 20551, 20206, 20400, 20804, 21911, 22864, 22010, 20933, 20173, 20059, 21233, 21651, 22336, 22609, 23121, 22749, 22388, 22728, 26561, 27107, 29304, 24449, 36625, 11837, 12431, 32358, 18405, 15362, 683, 9547, 7855, 3459, 4908, 3653, 3751, 3655, 3626, 3799, 3442, 4155, 1836, 0, 228, 0, 65, 0, 15, 0, 3, 0, 5, 0, 215, 1215, 629, 0, 79, 0, 23, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 169, 0, 609, 0, 5043, 11506, 8686, 9353, 18424, 25092, 20603, 19614, 20746, 20246, 19514, 19842, 20585, 20759, 21399, 21606, 21527, 22525, 23007, 22724, 22561, 22456, 22291, 22326, 22314, 22354, 22236, 22410, 23382, 29925, 13897, 584, 7040, 7111, 6142, 5435, 6679, 5612, 5473, 5626, 5895, 2697, 0, 3110, 2710, 0, 394, 0, 114, 0, 23, 0, 0, 0, 12, 0, 70, 0, 251, 0, 1636, 1768, 504, 1498, 148, 23, 0, 3, 2, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 108, 0, 402, 0, 3263, 8287, 10921, 9534, 6251, 7205, 6987, 6627, 7691, 5334, 13221, 20697, 17091, 17659, 17872, 18035, 18690, 20588, 21601, 22497, 22831, 22892, 22770, 21396, 24754, 27469, 26540, 26170, 25993, 27972, 27355, 28766, 22716, 18932, 18591, 16769, 10491, 2246, 9827, 17831, 6687, 0, 722, 0, 212, 0, 51, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 194, 0, 652, 0, 5627, 14169, 10684, 15431, 20151, 26367, 31605, 31006, 29323, 26233, 25747, 25253, 24053, 21830, 20001, 19160, 17990, 17059, 16860, 17005, 17730, 20941, 20439, 20182, 21522, 23296, 9112, 0, 1192, 0, 402, 113, 7, 836, 763, 0, 114, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 69, 0, 246, 0, 2371, 6117, 3086, 5315, 20523, 29512, 28601, 28644, 28370, 28769, 28794, 28743, 29059, 28334, 29728, 27135, 32319, 15339, 0, 4410, 2687, 4694, 3774, 4118, 4432, 4055, 4762, 5849, 5067, 4224, 4450, 5807, 2915, 5979, 0, 16849, 28077, 13592, 12872, 11895, 20924, 21528, 22641, 22497, 24155, 12068, 1363, 4509, 2081, 2996, 1196, 0, 149, 0, 49, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 107, 0, 919, 2625, 4899, 6479, 11027, 15231, 10757, 16384, 17393, 22640, 32650, 31597, 29999, 26910, 28129, 29184, 27051, 29538, 28389, 35848, 16677, 0, 2945, 270, 2264, 1849, 1462, 407, 1449, 3044, 5192, 5580, 6206, 4413, 6772, 0, 17345, 31507, 20871, 23916, 21883, 23331, 21930, 24025, 17697, 10649, 8591, 5628, 2663, 0, 343, 0, 68, 0, 11, 0, 0, 2, 0, 7, 0, 48, 48, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 48, 804, 9684, 17132, 14771, 12681, 12771, 17938, 19731, 19390, 20965, 20918, 22283, 23279, 22395, 22876, 24569, 24889, 25048, 24984, 25024, 24979, 25066, 24825, 24789, 23722, 25860, 25196, 28073, 25582, 28123, 22475, 4738, 6023, 6671, 5903, 5880, 5371, 6253, 2786, 0, 276, 0, 80, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 91, 0, 311, 0, 4518, 21651, 29986, 27232, 26287, 23426, 21601, 22474, 23258, 24759, 26650, 29201, 28551, 28183, 28551, 29274, 30618, 32194, 28870, 24254, 23381, 22823, 22908, 23958, 24346, 25773, 26804, 26395, 28795, 33680, 26341, 10955, 7256, 6709, 4229, 2396, 1626, 1422, 1405, 1423, 1393, 1463, 1329, 1601, 708, 0, 88, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 79, 0, 193, 0, 2924, 14305, 14056, 14012, 2957, 8019, 23883, 18971, 20401, 19822, 20120, 20267, 20059, 20218, 20811, 23727, 26347, 26377, 25262, 23965, 24027, 24174, 24087, 24217, 23997, 24347, 23724, 25495, 22633, 6170, 799, 3523, 13745, 24682, 16423, 6988, 4821, 3060, 1240, 1833, 630, 0, 57, 0, 20, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 14, 0, 60, 0, 413, 773, 1408, 826, 0, 113, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 227, 0, 795, 0, 6275, 13471, 10596, 11832, 11356, 11262, 11958, 10276, 15980, 21507, 19759, 20802, 21016, 21713, 21624, 22592, 23379, 23601, 23739, 22742, 22865, 22989, 22303, 22693, 21962, 22145, 21276, 23456, 25652, 27495, 15101, 5703, 9570, 7052, 6936, 7094, 6448, 5308, 4753, 4200, 3671, 1571, 54, 26, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 4, 0, 21, 0, 76, 0, 503, 503, 0, 76, 0, 21, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 157, 0, 448, 0, 4699, 13419, 716, 9243, 24830, 22401, 21476, 18851, 20266, 20151, 20048, 19616, 20129, 21983, 22394, 22076, 22625, 22831, 22464, 22018, 22242, 21769, 21172, 21287, 21222, 21467, 21834, 21887, 22047, 21666, 22409, 21025, 23809, 14420, 3114, 3945, 1652, 1924, 1048, 1937, 2709, 730, 0, 60, 0, 20, 0, 5, 0, 0, 0, 0, 8, 0, 49, 0, 179, 0, 2482, 6059, 7751, 8517, 7963, 5759, 1133, 0, 74, 0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 5, 0, 88, 0, 1656, 8902, 14112, 1047, 9360, 25781, 19403, 19148, 20036, 20332, 20259, 20315, 20199, 20451, 19900, 21727, 23545, 23047, 23339, 23535, 23585, 23510, 23609, 22828, 22595, 22597, 22585, 23567, 26831, 28001, 29582, 25642, 21217, 10095, 938, 6448, 7049, 7592, 11526, 16920, 17785, 16577, 20966, 10799, 0, 540, 0, 169, 0, 29, 0, 0, 0, 17, 0, 85, 0, 301, 0, 2340, 4790, 3198, 1306, 0, 167, 0, 42, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29729, 28756, 29021, 29343, 30109, 29864, 29423, 27373, 27753, 17661, 9426, 11332, 9064, 6439, 4361, 4827, 3119, 6387, 7639, 6223, 6971, 6350, 6710, 6393, 6799, 6141, 7409, 3277, 0, 407, 0, 116, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 154, 0, 533, 0, 4646, 12324, 11273, 11319, 11286, 11074, 11622, 10547, 12711, 5620, 0, 698, 0, 199, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 199, 200, 0, 32, 0, 0, 120, 0, 460, 0, 1583, 0, 12871, 29604, 30924, 29377, 37992, 12439, 11661, 38288, 26198, 29305, 27240, 27839, 26824, 27092, 27547, 27691, 27848, 27791, 27466, 26958, 27007, 27175, 27125, 26867, 27139, 27334, 27275, 27427, 27171, 27349, 27232, 27054, 27219, 27327, 27337, 27250, 27077, 26895, 26884, 26871, 26897, 26849, 26936, 26761, 27369, 28269, 28450, 28514, 28168, 28312, 28849, 28833, 28558, 27444, 25123, 9013, 0, 718, 0, 164, 0, 0, 264, 0, 3131, 8342, 8559, 11200, 6975, 5279, 3148, 0, 458, 0, 123, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 49, 449, 634, 1453, 3341, 8059, 11616, 11241, 12403, 12264, 12519, 13705, 12100, 9592, 8656, 8837, 8839, 8689, 9062, 8007, 8427, 9288, 9248, 6665, 1094, 0, 43, 0, 17, 0, 10, 0, 17, 0, 182, 572, 215, 0, 42, 0, 102, 0, 348, 0, 2802, 6309, 5676, 5441, 8896, 17607, 22605, 24389, 24662, 24549, 24327, 24527, 24536, 24866, 25144, 25219, 24849, 25715, 23906, 28525, 28250, 34547, 17061, 0, 4842, 0, 15828, 33760, 28054, 29080, 26896, 29104, 28852, 29727, 29780, 30184, 29896, 29055, 28604, 27906, 26215, 25357, 24622, 24492, 22413, 20564, 20555, 20388, 21069, 22742, 23853, 23174, 22578, 21262, 18240, 15194, 5986, 317, 1920, 1104, 1598, 1240, 1620, 688, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 97, 0, 788, 1770, 1488, 1597, 1597, 1488, 1770, 763, 0, 0, 180, 0, 815, 0, 7184, 19632, 23131, 28363, 30291, 31653, 31480, 31327, 31073, 30188, 28701, 28755, 29537, 30297, 29666, 24109, 6843, 0, 652, 0, 126, 0, 0, 387, 0, 3492, 10080, 17192, 25593, 26916, 28239, 28799, 28649, 28748, 28657, 28757, 28596, 29041, 29288, 29100, 29251, 28884, 29315, 27386, 30344, 24922, 36642, 12715, 11229, 35291, 26052, 25004, 17195, 20176, 18045, 17535, 17110, 16819, 16744, 15639, 13810, 13981, 12987, 12027, 11634, 13314, 17201, 20289, 18056, 10091, 0, 21398, 20210, 0, 3028, 0, 862, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 98, 0, 860, 3663, 12413, 19618, 21657, 23747, 25181, 29501, 26490, 34020, 15395, 0, 3124, 474, 2480, 1666, 2125, 2079, 1655, 2143, 177, 2689, 0, 14922, 33484, 27753, 30665, 28562, 28927, 28694, 28846, 28728, 29147, 29912, 29825, 29906, 29877, 30477, 30977, 30853, 30866, 30947, 30742, 31186, 29700, 28311, 29043, 28972, 28897, 29420, 28322, 27350, 27860, 27950, 28367, 28566, 28565, 29118, 29502, 29510, 29114, 26687, 25628, 23871, 22411, 18998, 15932, 17227, 13943, 3746, 0, 365, 0, 206, 0, 1000, 2973, 5729, 6937, 8708, 6826, 4477, 5936, 5318, 5624, 5492, 5502, 5634, 4718, 1237, 0, 110, 0, 32, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 63, 0, 217, 0, 3282, 16384, 24411, 26399, 27429, 27619, 28452, 28576, 28789, 28482, 29244, 28456, 30417, 26234, 35154, 11226, 11131, 35139, 26550, 30665, 27823, 28655, 28226, 28069, 28043, 27924, 27671, 27087, 26727, 26555, 25993, 25995, 25918, 25756, 25848, 25735, 25911, 25583, 26667, 27935, 27699, 28624, 28757, 29185, 29460, 29372, 29122, 28990, 29295, 29199, 29462, 28562, 28209, 28308, 28284, 28496, 27945, 26225, 25554, 25371, 24331, 19696, 19266, 7730, 0, 935, 0, 311, 0, 219, 0, 1337, 2965, 2562, 3140, 3477, 3217, 2823, 2880, 2964, 2720, 3257, 1446, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 181, 0, 644, 0, 5590, 15414, 18416, 21927, 22115, 23000, 24139, 24678, 26925, 28990, 29354, 30287, 30529, 31270, 32736, 30316, 28103, 28985, 28669, 28927, 28812, 28898, 29066, 29242, 29244, 29119, 29017, 29002, 29109, 29060, 29175, 29091, 29070, 29080, 29416, 29604, 29615, 29759, 29691, 29741, 29677, 29798, 29551, 30079, 28237, 22424, 6732, 0, 688, 0, 195, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 105, 0, 370, 0, 2940, 6755, 6916, 9300, 8598, 10484, 11568, 10073, 10178, 8487, 6650, 7166, 4528, 2479, 3100, 2730, 3041, 2677, 3275, 1438, 0, 179, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 61, 0, 294, 0, 1019, 0, 8470, 19456, 15891, 19699, 27043, 26961, 34882, 17080, 0, 4858, 0, 16487, 33604, 27260, 30332, 28353, 29267, 28868, 29213, 29250, 29259, 29179, 28921, 29078, 29193, 29152, 29192, 29134, 29232, 29046, 29598, 29849, 29653, 29836, 29886, 29789, 29651, 30125, 29869, 29617, 28734, 27427, 24015, 25256, 14999, 773, 261, 0, 92, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 86, 0, 310, 0, 2330, 4340, 3446, 3700, 3914, 1910, 0, 246, 0, 66, 0, 0, 63, 0, 353, 0, 1250, 0, 9978, 22754, 22543, 27475, 26185, 26737, 26772, 27588, 27786, 27843, 27737, 27664, 27731, 28081, 28284, 28306, 27896, 27048, 26932, 25972, 25259, 25477, 25342, 25465, 25298, 25601, 24666, 23170, 20579, 22430, 26477, 27644, 28501, 28471, 28440, 28706, 28207, 29436, 26860, 32802, 14354, 0, 3843, 1917, 2013, 4528, 0, 16727, 36685, 30362, 32253, 29576, 30273, 29576, 28382, 23000, 19920, 17664, 12005, 10252, 10627, 10158, 9609, 9073, 9185, 8922, 9402, 8527, 10275, 4546, 0, 564, 0, 161, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 134, 0, 521, 0, 7059, 23692, 28677, 30816, 29245, 36487, 16512, 0, 4430, 1399, 3171, 2226, 2136, 1707, 1881, 1879, 2312, 2663, 2873, 2916, 3086, 3002, 3038, 3088, 2942, 2827, 2961, 3092, 2779, 2965, 2902, 3214, 4256, 4613, 4466, 4717, 4184, 5250, 3232, 7135, 0, 14695, 32988, 26711, 30097, 28528, 29147, 28531, 28844, 29161, 29286, 28761, 30004, 28750, 28815, 19800, 3371, 0, 149, 0, 47, 0, 5, 0, 0, 68, 0, 239, 0, 2139, 6099, 7060, 7983, 8212, 8006, 8398, 8053, 7153, 7533, 7188, 7647, 6899, 8333, 3683, 0, 457, 0, 130, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2607, 2603, 2628, 2569, 2733, 2595, 2206, 2342, 2401, 1956, 1903, 2367, 2721, 2677, 2807, 2675, 2664, 1122, 0, 264, 0, 1111, 2469, 2648, 2983, 3133, 1637, 0, 1595, 1326, 0, 191, 0, 59, 0, 27, 0, 52, 0, 462, 1199, 809, 613, 705, 575, 799, 362, 1792, 3362, 3154, 3294, 2794, 2730, 2959, 2728, 3167, 3662, 3459, 3569, 3536, 3573, 3634, 3644, 3658, 3579, 3514, 3486, 3554, 3510, 3727, 3335, 3145, 1245, 0, 149, 0, 42, 0, 8, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1285, 2965, 2562, 2868, 2825, 3209, 3370, 3459, 3301, 3306, 2863, 2350, 2397, 2337, 2322, 2327, 2576, 2591, 2584, 2690, 2645, 3075, 3563, 3646, 3751, 3739, 3663, 3749, 3920, 3879, 3913, 4017, 3943, 3919, 3406, 3743, 1539, 0, 185, 0, 57, 0, 33, 0, 77, 0, 699, 2015, 2095, 2642, 2848, 2892, 2953, 3145, 3297, 3609, 3911, 3813, 3824, 3669, 3908, 3479, 2772, 2703, 2764, 2793, 2432, 3042, 3115, 2604, 2838, 2847, 3127, 2943, 3608, 4324, 3625, 3641, 3807, 3733, 3743, 3834, 3976, 3925, 3959, 3927, 3967, 3907, 4008, 3547, 2777, 3064, 994, 0, 0, 1423, 3447, 2926, 3416, 3358, 3478, 3283, 3430, 3599, 3668, 3843, 3766, 3720, 3149, 2812, 2975, 2935, 2870, 2950, 2861, 2872, 3102, 3003, 2992, 2901, 2927, 2895, 2841, 2861, 2850, 2955, 2962, 2955, 2976, 2933, 3015, 2850, 3389, 3918, 3746, 3861, 3996, 3990, 3979, 3832, 3529, 3766, 3722, 3507, 3274, 3164, 3274, 3391, 3493, 3466, 3450, 3387, 3551, 3630, 3747, 3890, 4122, 3965, 3821, 3441, 2928, 2930, 2705, 2616, 2702, 2742, 2715, 2850, 2728, 2730, 2849, 2807, 2829, 2818, 2822, 2823, 2826, 2891, 2891, 3252, 3685, 3601, 3812, 4042, 3996, 4113, 4198, 4253, 4290, 4082, 4147, 4156, 3827, 4136, 3845, 3307, 3282, 3287, 3437, 3434, 3410, 3289, 3320, 3279, 3532, 3670, 3673, 3894, 3721, 3713, 3101, 2719, 2902, 2689, 2656, 2650, 2661, 2643, 2677, 2608, 2838, 3095, 3111, 3125, 2975, 2869, 2700, 2676, 2797, 2596, 2995, 3471, 3481, 3466, 3472, 3755, 3746, 4134, 4552, 4617, 4603, 4528, 4531, 4538, 4169, 3749, 3590, 3277, 3268, 3285, 3134, 3157, 3377, 3340, 3264, 3413, 3301, 3450, 3619, 3576, 3581, 3610, 3536, 3695, 3165, 2649, 2928, 2952, 3180, 3119, 3111, 3174, 2888, 2862, 2932, 2823, 2864, 2804, 3206, 3626, 3560, 3600, 3713, 3672, 3748, 3837, 4291, 4683, 4653, 4774, 4883, 4740, 4700, 4885, 5380, 2045, 0, 290, 0, 756, 2622, 2718, 2278, 2407, 2365, 2350, 2431, 2234, 2895, 3500, 3467, 3446, 3447, 3647, 3593, 3175, 2997, 3301, 3184, 3157, 3320, 3198, 2691, 2536, 2610, 2418, 2361, 2750, 2747, 3149, 3461, 3451, 3564, 3548, 3800, 4020, 4158, 4504, 4849, 4687, 4894, 4166, 3446, 3532, 3541, 3850, 3828, 3897, 3775, 3999, 3583, 4412, 1830, 41, 598, 0, 0, 947, 2332, 1968, 2535, 2698, 2807, 2958, 3171, 3322, 3199, 3096, 3198, 2794, 2611, 2813, 2776, 2347, 1898, 1901, 2134, 2126, 2084, 2933, 2866, 2888, 3471, 3461, 3613, 3825, 4131, 4195, 4327, 3985, 3692, 3772, 3744, 3738, 3781, 3682, 4025, 4386, 3910, 4106, 3937, 4670, 1999, 0, 239, 0, 361, 808, 205, 482, 1898, 1875, 2311, 2894, 2946, 3043, 3215, 3393, 3523, 3572, 3459, 3339, 2995, 3055, 1274, 0, 767, 1422, 1478, 1894, 2663, 3082, 3007, 3337, 3503, 3459, 3485, 3461, 3492, 3440, 3573, 3593, 3728, 4011, 4047, 4270, 4041, 3832, 4474, 4037, 4667, 2051, 0, 255, 0, 73, 0, 14, 0, 3, 0, 13, 0, 219, 1263, 2507, 2984, 3053, 3159, 3215, 3334, 3269, 3369, 3078, 2862, 1212, 0, 907, 1695, 1482, 1623, 1477, 1681, 1317, 2487, 3844, 3758, 3918, 3700, 3683, 3446, 3580, 3842, 3840, 3897, 4077, 3828, 3718, 4283, 4141, 4540, 1782, 0, 210, 0, 60, 0, 11, 0, 0, 7, 0, 30, 0, 239, 707, 1827, 2918, 3003, 3113, 3176, 3358, 3414, 3410, 3395, 3432, 3355, 3514, 2998, 2459, 2374, 2762, 3302, 3082, 3322, 3634, 3645, 3789, 3856, 3449, 3671, 3451, 3731, 4101, 3861, 4196, 4136, 4151, 4298, 3821, 3647, 1364, 0, 158, 0, 45, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 57, 0, 198, 0, 1686, 4066, 2623, 1909, 2272, 1094, 0, 958, 2602, 805, 467, 2357, 2648, 2860, 3129, 3519, 3621, 3925, 3868, 3623, 1226, 0, 134, 0, 38, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 43, 0, 151, 0, 1261, 3067, 2818, 3081, 3277, 3727, 3720, 3753, 3682, 3550, 2851, 2622, 3014, 2730, 2714, 2732, 2528, 1975, 1991, 2294, 2362, 2488, 2958, 3456, 3499, 3642, 3758, 3739, 3526, 1189, 0, 129, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 158, 0, 1309, 3083, 2367, 2857, 3328, 3503, 3485, 3527, 3674, 2519, 2170, 2806, 2438, 2502, 2931, 2804, 2836, 2952, 2985, 2783, 2548, 2848, 2134, 2085, 2400, 2392, 2706, 2688, 3101, 3333, 3467, 3700, 3724, 3817, 3699, 3902, 3536, 4262, 1885, 0, 234, 0, 62, 0, 0, 38, 0, 157, 0, 1291, 3082, 2892, 3351, 3233, 3409, 3391, 3439, 3183, 2353, 2047, 2147, 2106, 2471, 2617, 2601, 2867, 2904, 2945, 2904, 2999, 2993, 3037, 3100, 3113, 3177, 3157, 3190, 3172, 3191, 3163, 3217, 3105, 3458, 3711, 3875, 3631, 4087, 1743, 0, 213, 0, 60, 0, 23, 0, 55, 0, 198, 0, 1535, 3184, 2688, 3264, 3338, 3279, 3075, 3388, 3417, 806, 746, 2671, 2388, 2739, 2891, 3131, 3090, 3141, 3205, 3202, 3278, 3305, 3300, 3291, 3317, 3263, 3372, 3062, 2957, 2587, 2304, 2554, 2654, 2655, 3131, 3661, 3410, 3606, 3396, 3877, 1569, 0, 187, 0, 60, 0, 42, 0, 112, 0, 928, 2347, 2663, 3253, 3125, 3577, 3298, 3287, 3174, 2680, 2426, 2160, 2705, 2798, 2667, 2680, 2664, 2679, 2664, 2684, 2646, 2802, 3136, 2995, 2962, 3050, 3042, 3091, 2938, 2810, 2708, 2718, 2749, 2786, 2771, 2844, 2873, 3252, 3614, 3516, 3579, 3429, 3444, 2867, 2792, 1143, 0, 112, 0, 0, 155, 0, 1446, 3469, 3085, 3451, 3339, 3584, 3369, 3097, 3229, 3077, 3308, 2915, 3660, 1402, 435, 2659, 369, 867, 2333, 1965, 2349, 2473, 2462, 2161, 1735, 2102, 883, 0, 66, 15, 0, 698, 2162, 2158, 2713, 3194, 3264, 3542, 3490, 3727, 3390, 2665, 894, 0, 99, 0, 27, 0, 5, 0, 0, 9, 0, 39, 0, 120, 0, 1186, 3394, 1121, 0, 0, 445, 1575, 1813, 2313, 2622, 2539, 2648, 2853, 2764, 2505, 2510, 2230, 2159, 868, 0, 93, 0, 0, 276, 1447, 1971, 2544, 3068, 3161, 3364, 3536, 3491, 3645, 3341, 4500, 2102, 0, 265, 0, 76, 0, 12, 0, 0, 18, 0, 65, 0, 656, 2240, 2733, 2464, 2465, 2800, 2468, 2351, 768, 0, 0, 742, 2480, 2472, 2438, 2234, 2817, 1208, 0, 153, 0, 66, 0, 92, 0, 725, 1943, 2097, 2604, 3124, 3496, 3423, 3426, 3580, 3619, 3653, 3560, 3745, 3398, 4093, 1811, 0, 225, 0, 64, 0, 10, 0, 0, 35, 0, 133, 0, 857, 967, 1037, 2248, 2152, 2532, 2135, 2653, 1100, 0, 90, 10, 0, 536, 564, 0, 76, 0, 0, 34, 0, 405, 1063, 901, 1713, 2244, 2092, 2178, 2112, 2181, 2077, 2454, 3322, 3426, 3569, 3555, 4068, 1647, 0, 196, 0, 56, 0, 11, 0, 0, 0, 0, 0, 0, 0, 3, 0, 8, 0, 15, 0, 424, 2216, 1116, 0, 140, 0, 41, 0, 9, 0, 0, 0, 10, 0, 47, 0, 160, 0, 1413, 3532, 2204, 2589, 4061, 3174, 3091, 3816, 3322, 3472, 3740, 3682, 3620, 2885, 3672, 1737, 0, 221, 0, 63, 0, 12, 0, 0, 0, 3, 0, 13, 0, 46, 0, 427, 1188, 1080, 1652, 2702, 2678, 2118, 2012, 2045, 1989, 2092, 1903, 2278, 1029, 0, 187, 0, 673, 2148, 2633, 2571, 3284, 1190, 0, 0, 1661, 3948, 3076, 3473, 3550, 3427, 3819, 1552, 0, 184, 0, 53, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 93, 0, 787, 2019, 1704, 2587, 1112, 0, 79, 31, 0, 1002, 3045, 2246, 1954, 821, 0, 104, 0, 30, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 0, 42, 0, 554, 2079, 890, 0, 103, 0, 31, 0, 7, 0, 0, 6, 0, 24, 0, 74, 0, 778, 2400, 889, 0, 94, 0, 29, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 55, 0, 895, 1603, 389, 0, 27, 0, 9, 0, 3, 0, 0, 0, 0, 0, 2, 0, 5, 0, 12, 0, 288, 1449, 718, 0, 89, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 25, 0, 90, 0, 595, 595, 0, 90, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 198, 198, 0, 30, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 19, 0, 68, 0, 450, 450, 0, 68, 0, 19, 0, 3, 0, 0, 0, 0, 0, 1, 0, 5, 0, 19, 0, 125, 125, 0, 19, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 68, 633, 1429, 2018, 2193, 2176, 2138, 2240, 2037, 2451, 1085, 0, 134, 0, 38, 0, 7, 0, 1, 0, 8, 0, 28, 0, 424, 321, 0, 46, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 44, 0, 147, 0, 1224, 2670, 631, 0, 40, 0, 15, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 47, 0, 175, 0, 1129, 962, 39, 1004, 2360, 3010, 2596, 2805, 692, 0, 56, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 60, 0, 218, 0, 1457, 1475, 0, 599, 1961, 1133, 0, 147, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 56, 0, 206, 0, 1345, 1250, 0, 0, 651, 815, 0, 126, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1545, 1610, 1540, 1582, 1739, 1395, 2115, 740, 3287, 0, 14847, 31206, 25333, 28322, 26995, 26416, 27153, 24572, 24692, 10264, 0, 1048, 0, 301, 0, 59, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 6, 0, 86, 338, 214, 277, 251, 66, 132, 97, 117, 104, 115, 85, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 883, 0, 3138, 0, 20590, 20829, 0, 4379, 0, 2528, 1622, 2417, 2410, 2739, 3011, 3195, 2770, 2929, 3393, 3468, 3258, 3103, 3078, 2897, 2915, 2764, 2726, 2823, 2505, 2027, 1547, 1459, 1358, 1269, 1416, 1452, 1526, 1480, 1541, 1439, 1621, 1260, 2459, 3790, 3566, 3594, 3562, 3830, 3453, 3247, 3190, 3149, 3104, 2694, 2150, 634, 0, 64, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 30, 551, 1092, 1456, 1663, 1623, 1676, 1587, 1798, 1898, 1799, 1453, 1957, 644, 2210, 281, 7254, 16774, 15160, 17118, 19362, 21795, 22140, 21917, 23356, 24622, 23248, 22432, 23053, 20738, 24381, 10669, 0, 1983, 110, 1082, 639, 960, 827, 847, 901, 786, 1003, 566, 2021, 3544, 2950, 3484, 3801, 4065, 4148, 4260, 4227, 4182, 4219, 4130, 3927, 3861, 4049, 3818, 3635, 3543, 3330, 2873, 2184, 1656, 523, 0, 55, 0, 15, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 276, 0, 984, 0, 9449, 20790, 21221, 23631, 23583, 25941, 25032, 25743, 25783, 26446, 26853, 27422, 27371, 26713, 27220, 26444, 27800, 25349, 30207, 14310, 0, 3117, 688, 3432, 3786, 4028, 4341, 4403, 4496, 4355, 4151, 4178, 4107, 4127, 4211, 4169, 4263, 4387, 4188, 4417, 4298, 4450, 4557, 4314, 4482, 4498, 4532, 4234, 4150, 4002, 4104, 3705, 3688, 1507, 0, 182, 0, 51, 0, 10, 0, 39, 0, 195, 0, 689, 0, 5565, 13113, 11388, 12682, 12055, 14342, 5546, 0, 653, 0, 193, 0, 54, 0, 170, 708, 1011, 1091, 1075, 1203, 1281, 1410, 1079, 748, 312, 0, 39, 0, 10, 0, 1, 0, 0, 0, 12, 0, 62, 0, 219, 0, 1793, 4282, 4181, 4679, 4501, 4836, 4906, 4797, 4794, 4585, 4060, 4436, 3718, 2846, 3159, 2734, 3377, 4525, 4663, 4997, 4950, 4613, 4682, 4317, 2410, 1258, 1442, 1348, 1429, 1537, 1480, 1593, 1682, 1813, 1768, 2458, 4236, 4767, 4660, 4700, 4689, 4676, 4727, 4500, 4064, 4164, 4071, 3771, 3344, 2968, 1763, 235, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 887, 0, 3151, 0, 20641, 20627, 0, 3857, 0, 1822, 533, 1124, 253, 0, 6, 32, 0, 245, 0, 884, 0, 7520, 19357, 20143, 22759, 24573, 26205, 26960, 26828, 27012, 23850, 25824, 11483, 0, 2509, 575, 1731, 1088, 1475, 1381, 1997, 2724, 3258, 3551, 3733, 4461, 4767, 4837, 4876, 5043, 5114, 5163, 5199, 5152, 5240, 5287, 5497, 5608, 5570, 5602, 5560, 5636, 5358, 4787, 4646, 4606, 4628, 4438, 4300, 3912, 3562, 1260, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 194, 0, 910, 0, 7333, 23432, 30566, 29528, 36790, 16379, 0, 2887, 314, 2322, 1942, 2069, 1527, 1895, 1077, 1916, 340, 2954, 0, 16469, 36143, 29004, 33121, 29262, 30892, 13262, 0, 3764, 2046, 3193, 2549, 2995, 3007, 3056, 3059, 3053, 3062, 3045, 3080, 2953, 2727, 2643, 2935, 3263, 3515, 3853, 4038, 4192, 4104, 4018, 4104, 4195, 3986, 3609, 1193, 0, 128, 0, 37, 0, 0, 47, 0, 252, 0, 875, 0, 7329, 17960, 15543, 16260, 15845, 15557, 15066, 15214, 15368, 14658, 13946, 14314, 13849, 14609, 13266, 15907, 7366, 0, 2657, 1697, 2230, 1674, 1894, 1771, 2020, 2169, 919, 304, 687, 112, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 1, 0, 4, 0, 137, 880, 1452, 1891, 2471, 2694, 2803, 2933, 3151, 3227, 3192, 3202, 3205, 3188, 3226, 3147, 3385, 3547, 3791, 4009, 3985, 4399, 4453, 3806, 3213, 3444, 3379, 3379, 2237, 975, 892, 1090, 1345, 2080, 3193, 3645, 4219, 4647, 4602, 4556, 4821, 4842, 4778, 4832, 4915, 4977, 4872, 4726, 4708, 4767, 4695, 4500, 4626, 4113, 3682, 3819, 3733, 3813, 3708, 3894, 3292, 2529, 2209, 1746, 606, 0, 67, 0, 18, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 92, 220, 163, 224, 131, 291, 0, 1010, 2165, 2044, 2029, 1710, 1740, 1977, 2078, 2117, 2026, 1882, 2068, 2401, 2544, 2596, 2576, 2599, 2541, 2431, 2662, 2388, 2322, 1976, 1620, 1690, 548, 0, 87, 0, 339, 1126, 1710, 2197, 2538, 2856, 3037, 3215, 3267, 3216, 3271, 3176, 3347, 3034, 3657, 1617, 0, 200, 0, 57, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 27, 0, 100, 0, 943, 2434, 2806, 3212, 3539, 2237, 857, 0, 1387, 0, 9904, 25243, 26922, 29474, 28436, 29034, 28601, 29074, 28318, 30618, 32815, 31923, 32079, 30119, 28452, 10519, 0, 2347, 581, 2176, 3275, 4210, 4440, 4368, 4328, 4374, 4241, 4064, 4087, 4226, 4334, 4421, 4479, 4502, 4366, 3977, 4012, 4185, 4151, 4153, 4165, 4164, 4036, 3890, 3804, 3724, 3657, 3632, 3678, 3580, 3769, 3419, 4119, 1822, 0, 226, 0, 64, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 13, 0, 44, 0, 465, 1638, 1914, 1984, 2163, 2288, 2618, 2560, 2696, 3017, 2815, 2858, 3051, 3084, 2901, 2907, 2822, 2751, 2778, 2715, 2941, 3138, 3166, 3163, 3166, 3161, 3172, 3145, 3254, 3367, 2820, 1793, 1342, 476, 0, 54, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 5, 1, 348, 1292, 584, 880, 0, 14875, 26450, 28530, 29079, 35789, 16866, 0, 3612, 541, 2147, 1040, 2028, 981, 1755, 0, 2375, 0, 16422, 36997, 30212, 33790, 27587, 30916, 13334, 0, 2196, 0, 1112, 295, 868, 243, 1921, 3709, 3310, 3494, 3393, 3664, 3595, 3606, 3785, 3733, 3655, 3610, 3519, 3375, 3378, 3335, 3092, 2921, 2241, 1865, 713, 0, 84, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 320, 0, 1113, 0, 8993, 20381, 16893, 18804, 15448, 4733, 0, 474, 0, 130, 0, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 64, 0, 307, 0, 1061, 0, 9357, 25538, 25071, 28260, 29472, 30450, 31537, 31538, 31427, 31296, 31309, 31326, 31316, 31317, 30782, 27769, 28017, 11117, 0, 2517, 613, 2176, 2609, 3051, 3338, 2988, 2789, 2857, 2570, 2643, 2817, 2884, 2997, 3076, 3228, 3276, 3363, 3520, 3665, 3598, 3506, 3413, 3277, 2570, 1996, 2054, 653, 0, 66, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 106, 0, 528, 0, 1857, 0, 14949, 34024, 29594, 32311, 30364, 30439, 28447, 28238, 27533, 28158, 27521, 25961, 8989, 0, 947, 0, 273, 0, 56, 0, 0, 0, 3, 0, 12, 0, 100, 91, 0, 13, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 0, 382, 0, 1348, 0, 10818, 25212, 22403, 25700, 23018, 24812, 9333, 0, 1094, 0, 315, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 594, 1147, 1324, 1383, 1752, 1969, 1662, 1643, 1515, 1376, 1736, 1728, 1578, 1807, 1896, 1977, 1888, 1740, 1821, 2125, 2073, 2199, 1577, 1247, 646, 0, 88, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 170, 0, 884, 0, 3139, 0, 20588, 20803, 0, 4283, 0, 899, 0, 156, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 0, 381, 0, 1335, 0, 11405, 29672, 29548, 31572, 30832, 32072, 31696, 31622, 31520, 31059, 30098, 28744, 27053, 25534, 9092, 0, 1671, 318, 1245, 1003, 2198, 3164, 3449, 3575, 3783, 3898, 3722, 3728, 3747, 3678, 3589, 3544, 3596, 3497, 3683, 3340, 4024, 1780, 0, 221, 0, 63, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 0, 189, 0, 668, 0, 7176, 19797, 24363, 28340, 28320, 29325, 29095, 29193, 29219, 29074, 28868, 29107, 24437, 26692, 11632, 0, 1373, 0, 391, 0, 92, 0, 1, 0, 7, 0, 173, 996, 1382, 1268, 1354, 1250, 1410, 1113, 2061, 2974, 2697, 2961, 2809, 2846, 2778, 2664, 2663, 2625, 2367, 1471, 317, 0, 24, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 137, 892, 1267, 1409, 576, 0, 70, 0, 21, 0, 15, 31, 97, 76, 174, 289, 252, 272, 259, 271, 253, 310, 378, 342, 219, 221, 31, 481, 1351, 1760, 1787, 1525, 1551, 1608, 1928, 2037, 1828, 615, 0, 67, 0, 19, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28246, 28894, 29871, 29592, 29574, 29422, 29624, 27441, 27776, 20452, 13905, 15694, 15118, 14862, 16180, 10997, 5185, 6593, 6244, 5719, 4473, 4768, 4249, 3637, 1201, 0, 131, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 27, 0, 76, 0, 1045, 4082, 1791, 0, 210, 0, 64, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 27, 0, 236, 563, 167, 36, 0, 249, 0, 2575, 2065, 8893, 14152, 10732, 14941, 19266, 35918, 15401, 0, 0, 15068, 35811, 26264, 28102, 27291, 28438, 27744, 27343, 27792, 28040, 27600, 27876, 28106, 28191, 28051, 27923, 27661, 27250, 27296, 27494, 27518, 27515, 27523, 27503, 27545, 27462, 27692, 27720, 27756, 27829, 27679, 28034, 27380, 26856, 26947, 27029, 26350, 25574, 25801, 25524, 25074, 25217, 25264, 25477, 25112, 25887, 26912, 26924, 26964, 27742, 24910, 21806, 17309, 4172, 0, 141, 172, 0, 3568, 10602, 7899, 5391, 4665, 4521, 4922, 4815, 4774, 4976, 4532, 5453, 2414, 0, 299, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 175, 0, 603, 0, 5070, 12533, 10668, 11707, 10221, 8437, 8115, 6743, 4447, 3923, 3635, 3306, 3698, 3089, 4229, 1892, 0, 235, 0, 18, 124, 0, 828, 0, 3096, 0, 20038, 18344, 0, 0, 15591, 34302, 15989, 5663, 0, 2112, 0, 7361, 13744, 11780, 13012, 11897, 13315, 10895, 18454, 25809, 22714, 23684, 23777, 23952, 24757, 26195, 28344, 31317, 31123, 33057, 30236, 35857, 16787, 0, 4841, 0, 17460, 35506, 29324, 31337, 28965, 25574, 21656, 22461, 21893, 21412, 21213, 21221, 20966, 20315, 20761, 20786, 21510, 23620, 24270, 24441, 24252, 24349, 24250, 24424, 24089, 24764, 22997, 23134, 19941, 18097, 9821, 0, 500, 0, 144, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 77, 0, 274, 0, 1797, 1797, 0, 272, 0, 59, 0, 0, 139, 0, 893, 1814, 9215, 14822, 15087, 14131, 20620, 26071, 34214, 16688, 0, 5196, 2413, 4078, 3184, 3632, 3560, 3889, 3453, 4090, 2083, 5105, 0, 15741, 34314, 28587, 31467, 29899, 30801, 30170, 30886, 29484, 31361, 29775, 36313, 16115, 0, 2925, 0, 3298, 0, 16933, 36975, 28690, 31133, 27863, 36511, 15848, 0, 2600, 3078, 0, 16450, 36058, 27969, 30646, 25419, 20450, 17715, 16860, 16548, 15798, 15196, 15038, 14298, 12844, 12443, 12022, 11735, 11946, 11602, 12217, 11101, 13319, 6038, 0, 694, 0, 199, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 215, 0, 814, 0, 6711, 15926, 20215, 24401, 33673, 15273, 0, 5040, 2720, 4848, 4207, 4772, 4673, 4918, 4930, 4920, 4592, 5241, 3730, 5877, 397, 16740, 33251, 28153, 30801, 29572, 30213, 29961, 29958, 30186, 29286, 28206, 28281, 28102, 28048, 28005, 27869, 27679, 27852, 27967, 28085, 28408, 28714, 28502, 28486, 28804, 29026, 29185, 29508, 29038, 28078, 28131, 28096, 28039, 28266, 28465, 28941, 28449, 28195, 25860, 24513, 25143, 23726, 21721, 19309, 17543, 16966, 17103, 16899, 17191, 16643, 17678, 15754, 19571, 7755, 477, 6841, 7106, 6250, 2329, 3998, 4704, 4508, 5191, 3305, 1420, 1323, 0, 215, 0, 54, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 594, 0, 2120, 0, 13833, 13681, 0, 4649, 1905, 4205, 3449, 4043, 3978, 4044, 3972, 3913, 4015, 3716, 3680, 1486, 4150, 0, 14486, 31819, 25768, 28316, 26900, 27610, 27338, 27321, 27595, 26588, 25716, 25761, 25067, 25451, 26122, 26641, 26861, 27089, 27423, 27414, 27437, 27596, 27648, 28257, 28333, 28463, 28403, 29344, 29690, 29107, 28810, 29037, 28849, 28226, 28367, 28652, 28070, 29660, 30388, 26944, 26018, 26410, 24836, 21708, 16641, 12826, 8740, 6170, 6965, 6483, 6908, 6374, 7290, 4583, 2585, 2477, 2089, 3312, 3431, 2872, 507, 0, 26, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 37, 0, 128, 0, 1528, 5901, 7786, 7316, 8174, 6533, 13726, 25104, 26446, 25638, 26406, 27600, 29877, 28008, 35579, 16060, 0, 2657, 377, 912, 2278, 0, 15009, 33388, 27637, 30232, 28364, 29350, 28856, 28880, 28854, 28843, 28844, 28854, 28828, 28884, 28705, 28593, 28764, 28798, 28885, 28889, 28806, 28806, 28717, 28783, 28674, 28804, 28933, 28694, 28702, 28312, 27998, 27960, 27563, 27259, 27790, 26905, 27280, 25377, 25822, 10013, 0, 1176, 0, 336, 0, 82, 0, 66, 0, 232, 0, 1863, 4253, 3454, 3985, 3463, 4182, 2904, 6755, 9203, 7581, 8596, 8042, 2946, 0, 332, 0, 91, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 50, 0, 242, 0, 858, 0, 7428, 18935, 18860, 18928, 25402, 28492, 35530, 16766, 0, 3957, 2268, 2396, 4676, 0, 16819, 36721, 30534, 33797, 31748, 33419, 30374, 28115, 28892, 28349, 28433, 28356, 28539, 28460, 28554, 28498, 28676, 28720, 28789, 28770, 28919, 29035, 28959, 29080, 29082, 28882, 29052, 28859, 29239, 28740, 29585, 23774, 11079, 8811, 3615, 0, 443, 0, 127, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 38, 0, 596, 2862, 3569, 4378, 5144, 5204, 5547, 5845, 2859, 487, 510, 0, 184, 0, 446, 0, 1427, 0, 12578, 33110, 25484, 29240, 32131, 27171, 25208, 25750, 25971, 29455, 14299, 0, 14681, 28909, 25106, 27016, 25878, 26639, 25980, 27306, 28443, 27859, 27958, 27646, 27392, 26931, 26545, 26361, 26081, 26097, 25936, 25902, 25994, 25604, 25973, 27028, 28262, 28588, 28486, 28727, 28534, 28639, 28395, 28449, 28849, 28796, 29450, 29431, 30470, 31587, 31037, 29557, 28653, 29092, 28110, 27939, 28226, 27968, 28275, 27761, 28671, 27025, 30350, 18575, 883, 360, 0, 126, 0, 8, 0, 0, 0, 1, 0, 9, 0, 35, 0, 255, 438, 301, 405, 357, 651, 287, 0, 35, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 35, 0, 310, 664, 4701, 15695, 25697, 25097, 33753, 16064, 0, 5800, 3238, 4916, 4151, 4604, 4502, 4558, 4627, 4754, 4810, 4487, 4101, 4064, 3824, 3674, 3724, 3683, 3734, 3656, 3758, 3417, 2552, 3360, 1744, 3990, 0, 14621, 33679, 28495, 29029, 28226, 28397, 28187, 28183, 28058, 27964, 28360, 27461, 29968, 25904, 35197, 16137, 0, 0, 13592, 33184, 26652, 29648, 27899, 27628, 28767, 26800, 31598, 13596, 0, 1668, 0, 466, 0, 28, 92, 0, 489, 0, 3828, 8447, 8232, 6621, 2565, 1078, 0, 363, 154, 0, 16, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 334, 0, 3043, 9046, 10904, 11362, 11369, 11075, 10522, 11023, 11238, 12980, 14080, 14337, 14221, 11361, 10370, 5262, 1273, 1187, 0, 202, 0, 48, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 40, 0, 135, 0, 1452, 5426, 6281, 6820, 6495, 6989, 3874, 1616, 1966, 4374, 3583, 11795, 21859, 22676, 26326, 26248, 27645, 28550, 29040, 29282, 29825, 30524, 30934, 31210, 30944, 31399, 30583, 32173, 27234, 23740, 26296, 25422, 25836, 17379, 15588, 16929, 18046, 18335, 22502, 10920, 0, 1253, 0, 356, 0, 70, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 124, 0, 433, 0, 3355, 6787, 4482, 4978, 3994, 3017, 3011, 3108, 3524, 2556, 4445, 627, 12802, 22599, 17737, 13988, 9708, 8479, 3644, 2876, 2089, 1021, 0, 126, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 157, 0, 547, 0, 4559, 11109, 9241, 10012, 10816, 14745, 14750, 17001, 21839, 23405, 25547, 26805, 23183, 20108, 17384, 9655, 7137, 8336, 8999, 9404, 9305, 9160, 8756, 8874, 7914, 5492, 4540, 3845, 2799, 4100, 1954, 0, 246, 0, 71, 0, 14, 0, 0, 0, 0, 0, 4, 0, 20, 0, 69, 0, 623, 1714, 1487, 1635, 2017, 2053, 2062, 1766, 2356, 1318, 0, 818, 3589, 7071, 9258, 11015, 11563, 12002, 12462, 13058, 14415, 15391, 16222, 16701, 16209, 17277, 12771, 7798, 7152, 5203, 5464, 5338, 6735, 6192, 4857, 5358, 5001, 5377, 4844, 5818, 2633, 0, 1844, 2829, 2763, 2966, 3145, 3042, 3298, 2609, 2004, 1375, 0, 3520, 14640, 21091, 17331, 7914, 4444, 1938, 135, 2201, 1832, 2756, 1190, 0, 65, 0, 6, 17, 0, 105, 0, 1021, 3239, 4086, 4380, 4840, 5293, 5170, 5198, 5243, 5106, 5413, 4357, 2749, 939, 0, 88, 0, 0, 230, 345, 789, 1855, 1922, 2100, 2101, 2924, 4213, 2555, 314, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 232, 1813, 4228, 5072, 4808, 5066, 4696, 5312, 4138, 7957, 11701, 9716, 11454, 6017, 71, 184, 0, 66, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 52, 0, 188, 0, 1379, 2408, 1709, 1934, 2396, 3512, 3274, 2915, 3974, 4171, 4117, 2102, 0, 117, 0, 0, 440, 723, 2268, 4388, 4639, 4634, 3984, 1313, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 114, 0, 400, 0, 3278, 7799, 6982, 7941, 7847, 8725, 7721, 10850, 13581, 10742, 16475, 19671, 18221, 18858, 17800, 17377, 17592, 17616, 18744, 13171, 3615, 5519, 10141, 10675, 10292, 9694, 10115, 10573, 10441, 10512, 10464, 10503, 10507, 9661, 3423, 0, 949, 155, 28, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 5, 0, 51, 0, 235, 0, 1251, 467, 5487, 11977, 16407, 23321, 24567, 25379, 26023, 27241, 29481, 30340, 31314, 32582, 32075, 31723, 31235, 31451, 31249, 31528, 31060, 31973, 28890, 24602, 22450, 18579, 18230, 18450, 17682, 16721, 16504, 15009, 14405, 12995, 11334, 12249, 8707, 2686, 67, 29, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 36, 50, 1199, 1141, 2317, 3277, 3659, 4744, 4411, 4487, 4618, 4235, 5077, 2251, 0, 279, 0, 79, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 53, 0, 176, 0, 1489, 3578, 2147, 3157, 2676, 1540, 2159, 2861, 1143, 0, 0, 549, 0, 5292, 13149, 12478, 13024, 14064, 13246, 15033, 6674, 0, 828, 0, 220, 0, 0, 138, 144, 1014, 1773, 1530, 1445, 1017, 1077, 1261, 1301, 1311, 1277, 1344, 1219, 1469, 650, 0, 80, 0, 22, 0, 14, 0, 48, 0, 136, 0, 1730, 4515, 3202, 4617, 689, 5239, 15984, 14961, 16243, 21597, 25367, 26862, 27130, 26911, 26499, 25801, 23903, 20123, 18598, 18133, 18235, 19001, 19287, 17590, 16869, 15407, 13840, 14491, 13870, 14735, 13297, 16070, 7088, 0, 834, 0, 1440, 401, 0, 40, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 491, 663, 951, 2261, 2706, 4210, 5857, 6332, 5859, 5336, 5830, 5412, 5585, 5560, 5027, 4929, 4897, 4989, 4807, 5150, 4473, 6462, 6623, 3978, 3837, 4151, 3244, 3099, 3698, 4332, 4719, 1999, 284, 0, 10, 0, 0, 10, 0, 75, 99, 0, 100, 0, 314, 0, 2139, 2092, 0, 306, 0, 49, 28, 0, 582, 1310, 702, 1436, 2141, 2077, 2139, 2087, 2144, 2062, 2212, 1695, 923, 776, 208, 0, 18, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 3, 0, 18, 0, 62, 0, 697, 2686, 3483, 3738, 3773, 3916, 3724, 4063, 1641, 0, 192, 0, 55, 0, 11, 0, 0, 0, 0, 3, 0, 39, 0, 362, 1002, 2248, 1020, 5882, 9770, 7157, 5982, 4484, 4804, 4214, 3444, 3156, 2777, 2903, 3333, 2965, 2391, 1759, 1146, 266, 0, 22, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 34, 0, 134, 0, 1035, 2491, 4233, 3395, 2010, 4149, 7376, 11064, 14194, 15596, 16779, 18514, 18459, 18116, 20589, 20147, 19912, 19419, 19425, 21476, 21463, 21927, 19397, 18794, 17565, 16035, 14851, 14029, 14009, 13892, 13633, 14294, 12991, 15639, 6922, 0, 859, 0, 246, 0, 49, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 66, 0, 306, 0, 1393, 0, 8807, 17664, 15583, 18046, 17929, 18944, 19735, 19145, 21651, 24039, 23365, 23626, 23620, 23345, 24504, 25474, 24808, 25484, 23978, 21478, 19954, 21518, 19768, 20072, 24272, 21980, 25421, 14635, 3013, 6724, 2320, 0, 4300, 2645, 0, 335, 0, 103, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 0, 200, 0, 699, 0, 5784, 13786, 11895, 12375, 12035, 11809, 13333, 16274, 17591, 18410, 19097, 19828, 19180, 20742, 21556, 22010, 23512, 24802, 26468, 26578, 27274, 27319, 28312, 29597, 30434, 29912, 28814, 29426, 30870, 31911, 30947, 31923, 29374, 31156, 15825, 505, 0, 10251, 21294, 17713, 19801, 18092, 20107, 16936, 24077, 12977, 0, 1409, 0, 891, 3157, 2830, 7670, 11990, 5299, 2790, 3402, 3788, 6532, 5969, 12185, 19997, 22061, 23564, 20789, 13864, 10339, 11727, 11149, 11029, 10229, 10019, 5024, 2878, 3033, 647, 262, 0, 39, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 71, 0, 222, 0, 3075, 5438, 3651, 5225, 1233, 5469, 14403, 12904, 19277, 26289, 27818, 27676, 29292, 24888, 18275, 18702, 18030, 18515, 17978, 18779, 17398, 20112, 11300, 2963, 5837, 4248, 4567, 4151, 1645, 0, 183, 0, 52, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 62, 0, 235, 0, 1644, 2835, 3581, 2939, 879, 1306, 1617, 500, 2833, 0, 13962, 30476, 24480, 26823, 18833, 16324, 12337, 6939, 7873, 7286, 3158, 0, 320, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 304, 0, 1063, 0, 8491, 18564, 14432, 18957, 21814, 20053, 15305, 15139, 15610, 18483, 19317, 25280, 31834, 30884, 32395, 30464, 27880, 24504, 13318, 7993, 9081, 8272, 8144, 7817, 7180, 4849, 1870, 0, 61, 0, 17, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 47, 0, 193, 0, 1390, 3077, 7626, 13357, 15781, 17070, 17057, 16266, 15762, 16624, 15430, 13131, 13547, 15334, 14542, 15407, 8053, 2322, 4180, 3885, 4604, 4956, 5243, 5330, 5221, 5385, 5881, 5857, 5744, 5487, 4802, 3653, 1035, 0, 101, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 20, 0, 97, 0, 322, 0, 2888, 7922, 6826, 9563, 10197, 9007, 10012, 9728, 10888, 11126, 11108, 9760, 9438, 7117, 6605, 4905, 10697, 16934, 16955, 20941, 22128, 24583, 27293, 29918, 30316, 30763, 30894, 30987, 30716, 31269, 30215, 32357, 25090, 15415, 12293, 9336, 9772, 8502, 8153, 7323, 5495, 4174, 3493, 3246, 2885, 2773, 1254, 0, 158, 0, 43, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 158, 477, 1835, 962, 5167, 10071, 9790, 10475, 10133, 10348, 10180, 10365, 10025, 11620, 15569, 12009, 7850, 8291, 8947, 9660, 10035, 10370, 10594, 10116, 9106, 8011, 6747, 6896, 6583, 6086, 5749, 4872, 5738, 2423, 0, 294, 0, 84, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 75, 0, 370, 0, 1304, 0, 10915, 27192, 26155, 27785, 27515, 28944, 26540, 25427, 23119, 22610, 22659, 22991, 22004, 21243, 21987, 20817, 20475, 19753, 19761, 19555, 19298, 19225, 18757, 17821, 17634, 17476, 16628, 12636, 10868, 12694, 11325, 9619, 3188, 0, 349, 0, 101, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 130, 0, 450, 0, 3432, 6626, 4199, 6090, 5053, 1463, 0, 1085, 3127, 4107, 6660, 9248, 10110, 10665, 12122, 12112, 11790, 13148, 14061, 13581, 10033, 2729, 0, 259, 0, 73, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 104, 0, 346, 0, 3144, 8727, 6790, 8414, 9434, 8985, 6673, 5944, 3693, 6328, 13606, 17574, 20540, 21582, 19817, 16586, 11670, 7902, 8840, 8706, 8182, 9681, 4326, 0, 535, 0, 153, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 0, 92, 295, 322, 261, 577, 2804, 3816, 3801, 3398, 4336, 2331, 9263, 17683, 16775, 17817, 18013, 17019, 17538, 13146, 9150, 8924, 9811, 4513, 0, 567, 0, 156, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 149, 0, 531, 0, 4247, 10052, 10194, 7232, 716, 18, 0, 2, 85, 229, 0, 1441, 0, 5000, 0, 22866, 21195, 0, 11166, 9357, 11385, 9915, 7570, 6251, 5062, 3811, 4060, 1161, 0, 106, 0, 34, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 3, 0, 158, 659, 518, 802, 0, 4002, 10840, 12173, 13472, 14129, 15230, 15290, 15951, 16604, 17162, 16242, 13773, 13419, 7399, 1044, 519, 0, 97, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 13, 0, 27, 502, 4908, 5733, 6682, 11241, 8609, 1983, 0, 1012, 1835, 4558, 6486, 7988, 9383, 9858, 9896, 9755, 9875, 9794, 9893, 9733, 10015, 9454, 11339, 13539, 12872, 11888, 10826, 10515, 9829, 9399, 8741, 8069, 8280, 6749, 1748, 0, 153, 0, 44, 0, 10, 0, 0, 0, 0, 0, 0, 27, 0, 131, 0, 457, 0, 3718, 8442, 7106, 11287, 14954, 15435, 14596, 14421, 14348, 14575, 14107, 14989, 13209, 19237, 26504, 25589, 26607, 26873, 26905, 25026, 20788, 16907, 11798, 10093, 4166, 0, 510, 0, 141, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 54, 0, 179, 0, 1518, 3443, 853, 0, 107, 980, 1152, 1152, 1104, 3504, 5863, 12850, 17958, 18624, 20353, 21910, 21201, 18547, 17094, 16906, 9082, 1240, 1146, 0, 210, 0, 45, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 135, 0, 495, 0, 3968, 9704, 11533, 14497, 15527, 20109, 13547, 1840, 3892, 10457, 12599, 14259, 14268, 12075, 11592, 11620, 10962, 10941, 10853, 10624, 10818, 10498, 11071, 10032, 12093, 5349, 0, 664, 0, 190, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 0, 0, 998, 8574, 12382, 11983, 7243, 3557, 7770, 6567, 3095, 1068, 2105, 3101, 6367, 6434, 6657, 10555, 11470, 12138, 11916, 11994, 12007, 11909, 12136, 11346, 10353, 10435, 9936, 10101, 10110, 10256, 8925, 7043, 2406, 0, 269, 0, 75, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 103, 0, 383, 0, 2308, 1423, 2912, 17162, 23812, 18622, 15750, 17178, 16336, 16661, 16764, 17956, 19784, 20350, 19644, 19338, 19688, 19663, 19593, 19393, 19587, 18616, 18213, 18125, 18747, 19195, 20825, 23936, 24039, 24653, 22351, 21758, 25914, 13765, 5300, 7839, 5974, 6269, 5847, 6102, 5866, 6200, 5624, 6776, 2998, 0, 372, 0, 106, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 11, 0, 123, 0, 1601, 6978, 12347, 650, 10027, 25857, 21007, 22978, 18966, 18176, 18703, 19164, 19761, 19986, 20775, 20452, 20548, 20315, 20371, 20415, 20251, 20616, 19630, 19739, 19498, 23096, 26178, 23895, 24509, 24326, 22794, 23596, 18198, 8373, 6609, 6427, 3596, 3634, 5314, 4089, 3566, 3402, 4104, 1812, 0, 226, 0, 63, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 238, 0, 918, 0, 5252, 2498, 6425, 22731, 24618, 29132, 28631, 28834, 28303, 26767, 24731, 22992, 23478, 22946, 21913, 22224, 21424, 21162, 20737, 19403, 18648, 18012, 18000, 19325, 22164, 27330, 22537, 32040, 9984, 13514, 35347, 18312, 20200, 9352, 4033, 5241, 3536, 3162, 1587, 880, 1049, 996, 965, 1124, 507, 0, 62, 0, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 62, 0, 330, 0, 1214, 0, 8856, 15847, 15125, 19878, 23041, 29849, 27423, 27488, 27705, 27837, 27783, 27226, 26217, 26020, 26061, 25482, 24404, 22945, 21893, 22090, 22413, 22508, 22408, 22659, 22110, 23187, 21069, 26923, 29338, 34001, 19136, 0, 18838, 30940, 16098, 6393, 577, 2137, 1145, 2186, 3200, 3171, 3993, 1781, 0, 222, 0, 64, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 163, 0, 572, 0, 4576, 10499, 8445, 9925, 8305, 10682, 6316, 20010, 31544, 25606, 27506, 29682, 31232, 31145, 32612, 31845, 25906, 34077, 12508, 9292, 42985, 11874, 11336, 40276, 13711, 0, 1853, 5809, 1228, 18487, 32112, 20127, 24108, 20390, 20041, 7899, 0, 1763, 355, 1263, 1236, 633, 0, 71, 0, 20, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 59, 0, 243, 0, 2810, 11019, 15802, 14228, 22596, 31495, 30017, 31304, 29737, 27823, 26719, 23798, 22740, 22462, 23147, 23613, 21741, 22684, 23093, 21619, 20846, 21004, 21736, 23784, 27121, 30143, 32025, 32321, 32409, 32133, 32695, 31648, 33756, 26530, 17220, 18858, 18174, 17220, 6079, 0, 715, 0, 183, 0, 61, 0, 50, 173, 3196, 6139, 5163, 5331, 2104, 0, 252, 0, 74, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 170, 0, 570, 0, 4498, 9965, 6496, 4462, 0, 10199, 26596, 25575, 25851, 25572, 25599, 25831, 25280, 26425, 22593, 18187, 19053, 19319, 20826, 21054, 22437, 23416, 24707, 25691, 25866, 26035, 25668, 26438, 26836, 27976, 30771, 25417, 18190, 24557, 30348, 22503, 19835, 13430, 2571, 1973, 1566, 1462, 1089, 1024, 815, 945, 402, 0, 48, 0, 14, 0, 2, 0, 11, 0, 56, 0, 195, 0, 1430, 2257, 138, 55, 0, 17, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 66, 0, 247, 0, 2406, 6683, 5218, 5362, 18517, 27473, 25510, 26111, 25824, 25096, 23208, 22129, 21959, 21527, 21379, 21779, 22388, 22840, 22038, 20508, 20553, 21195, 21052, 21083, 21443, 22357, 22118, 21243, 21348, 24238, 28947, 25714, 34176, 15959, 0, 3347, 190, 1945, 919, 1609, 903, 2633, 4073, 4535, 5396, 4959, 5028, 5158, 4498, 5432, 2480, 0, 312, 0, 89, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 93, 0, 390, 0, 3396, 8763, 10301, 3318, 13042, 26704, 24360, 25742, 22309, 20832, 19916, 20905, 22966, 23355, 23246, 23411, 23109, 23698, 21916, 20999, 21780, 20707, 21081, 22231, 22948, 24999, 27478, 25773, 29679, 30304, 28564, 18893, 6662, 6381, 5633, 4565, 5600, 6389, 5519, 5380, 5731, 3051, 0, 3121, 2621, 0, 378, 0, 111, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 164, 0, 565, 0, 8181, 17371, 17280, 20274, 20943, 22339, 17010, 17514, 21048, 19002, 19848, 19286, 19710, 19936, 19189, 19581, 21066, 20873, 21402, 22512, 21587, 21766, 22677, 24051, 23404, 24967, 27391, 26345, 26988, 27027, 23931, 17978, 17256, 15878, 20413, 19041, 13483, 16161, 14576, 15987, 14205, 17283, 7613, 0, 947, 0, 271, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 101, 0, 272, 1204, 19114, 30790, 28445, 31701, 31060, 31477, 29462, 27346, 26707, 25682, 23358, 21785, 22419, 22407, 21608, 20333, 19994, 20022, 20086, 19932, 20237, 19613, 21847, 24828, 22900, 20984, 14410, 5703, 4367, 4108, 2049, 1407, 1559, 630, 0, 70, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 98, 0, 484, 0, 1692, 0, 13629, 30806, 25435, 28306, 26954, 26749, 23819, 25192, 22594, 36422, 13565, 9159, 39755, 12660, 307, 4633, 3382, 4200, 2700, 3718, 5088, 5252, 5418, 5928, 3322, 4943, 0, 18379, 35529, 24563, 23417, 13167, 15663, 22590, 22894, 23437, 22496, 21053, 18560, 19590, 18691, 19878, 17936, 21664, 9574, 0, 1190, 0, 340, 0, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 36, 0, 92, 0, 1587, 7474, 8865, 13647, 14767, 18503, 26740, 27791, 28150, 27295, 26007, 24349, 25777, 26528, 23625, 24451, 26679, 27742, 29230, 29425, 29187, 28822, 30354, 30292, 29319, 29645, 29907, 30291, 29202, 31467, 27146, 35589, 11898, 13240, 30052, 16101, 21101, 17715, 17994, 15801, 16276, 14389, 13238, 7436, 686, 149, 0, 30, 0, 0, 0, 0, 21, 0, 112, 0, 383, 0, 3059, 7060, 6115, 6586, 2008, 0, 204, 0, 65, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 148, 0, 510, 0, 4403, 11606, 10836, 9923, 6795, 3457, 2316, 2356, 2755, 1813, 3637, 0, 12357, 25946, 21802, 23185, 22186, 22714, 23417, 23559, 22981, 23130, 24025, 24106, 25609, 23941, 26813, 25513, 35209, 10729, 12530, 32553, 8778, 5918, 4817, 5232, 5812, 3001, 0, 172, 0, 57, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 0, 70, 0, 289, 0, 4343, 1039, 5822, 25135, 29328, 27920, 27461, 26108, 26594, 26155, 25789, 28994, 30452, 30854, 30958, 29860, 29106, 28717, 27577, 27048, 25614, 23688, 23712, 23069, 24143, 23698, 26265, 28836, 28297, 29148, 28647, 29154, 28394, 29710, 27328, 32078, 16305, 0, 2633, 740, 1047, 0, 156, 0, 20, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 135, 0, 452, 0, 3559, 8234, 5877, 4303, 0, 11415, 25706, 20810, 21797, 21062, 21210, 21067, 21194, 21004, 21352, 20618, 23150, 25852, 23212, 22202, 22217, 21608, 22946, 24646, 24947, 24741, 26457, 26829, 27728, 26875, 31961, 24530, 20178, 14460, 4831, 5914, 2347, 2880, 999, 1764, 588, 0, 67, 0, 21, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 63, 0, 149, 0, 1932, 6031, 0, 9689, 25658, 24349, 25284, 24304, 22858, 21413, 21531, 21322, 21425, 21612, 21327, 21520, 22482, 22875, 23515, 24602, 23558, 22862, 22958, 22576, 22668, 21787, 21340, 21883, 22646, 26695, 26545, 28256, 25572, 20477, 14556, 7371, 6657, 5287, 5683, 5707, 5294, 6319, 2806, 0, 348, 0, 99, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 138, 0, 422, 0, 3287, 5098, 0, 12843, 25796, 21912, 24048, 22880, 22277, 21543, 21161, 21566, 21760, 22647, 22769, 22862, 23278, 23145, 23189, 23209, 23115, 23326, 22660, 22160, 22387, 21440, 22276, 25050, 28927, 28746, 10574, 755, 5318, 5862, 14627, 9564, 766, 2411, 2491, 2697, 1602, 697, 0, 80, 0, 22, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 434, 0, 1511, 0, 12101, 26749, 20416, 22116, 20753, 21502, 21416, 21690, 22504, 24321, 24476, 24626, 25161, 25344, 25833, 24971, 24788, 24998, 24236, 23286, 23518, 23859, 23601, 23706, 25091, 25178, 29860, 27951, 7593, 0, 4175, 6763, 4398, 9564, 20845, 19074, 16561, 16844, 17060, 17225, 16775, 17656, 16015, 19290, 8537, 0, 1060, 0, 303, 0, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12897, 12922, 12828, 12700, 12579, 12047, 8762, 6707, 7162, 9372, 11591, 11988, 12687, 12979, 12712, 12348, 12245, 12263, 11826, 11485, 11408, 11042, 10456, 11230, 6334, 1250, 0, 5309, 13918, 13191, 13803, 13519, 13555, 13749, 13232, 15037, 16901, 16140, 16010, 15927, 15922, 15368, 13820, 11407, 12713, 17074, 18871, 17738, 16704, 17521, 14361, 11450, 12439, 11282, 14042, 6441, 0, 619, 0, 177, 0, 7, 34, 0, 173, 0, 1518, 4079, 3900, 5509, 5914, 7430, 10864, 11599, 11559, 11465, 11693, 11242, 12171, 9014, 5339, 5976, 5604, 5868, 5691, 5815, 5827, 5817, 5179, 5298, 5437, 2438, 1026, 499, 0, 312, 184, 343, 553, 774, 798, 415, 690, 1353, 1597, 2145, 2311, 2666, 2468, 2154, 1874, 3073, 3828, 3685, 4078, 4786, 2950, 1160, 1668, 1479, 1464, 1687, 1133, 2939, 4023, 3091, 3493, 3123, 3269, 3185, 3293, 3209, 3359, 3410, 3089, 2953, 2903, 3020, 3210, 4446, 3773, 2171, 2399, 2156, 1850, 2040, 2064, 2118, 2499, 2569, 2826, 2597, 2759, 5021, 6438, 6244, 6160, 6439, 6537, 6451, 6602, 6639, 6634, 6636, 6634, 6638, 6629, 6665, 6729, 6829, 6641, 6584, 6097, 6594, 5028, 3186, 3288, 2744, 3087, 2838, 2809, 3154, 2410, 2383, 2682, 2102, 2097, 2169, 3719, 3498, 3623, 1512, 116, 795, 0, 149, 0, 41, 0, 28, 0, 81, 0, 1075, 3418, 3909, 3815, 3907, 3761, 4016, 3520, 5127, 6717, 6291, 6487, 5950, 5672, 5689, 4385, 1068, 0, 89, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 9, 45, 559, 343, 0, 46, 0, 13, 0, 2, 0, 0, 11, 0, 58, 0, 204, 0, 1701, 4162, 3741, 4007, 3846, 3963, 3841, 4014, 3780, 4936, 3412, 216, 52, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 18, 0, 122, 122, 0, 13, 1, 0, 52, 0, 196, 0, 1594, 3557, 3186, 2668, 2833, 2426, 4412, 7655, 7814, 8177, 6661, 6548, 5749, 5976, 2616, 0, 415, 0, 412, 0, 2590, 5896, 4768, 5535, 4768, 5904, 2572, 0, 321, 0, 92, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 28, 0, 94, 0, 879, 2591, 2260, 3753, 4920, 5431, 3873, 2578, 3463, 3440, 3211, 4181, 3478, 7485, 11425, 9767, 10052, 9988, 10245, 10036, 9824, 9919, 11704, 12298, 12168, 11408, 10577, 10905, 10160, 9829, 9530, 10206, 10871, 10650, 10806, 10631, 10902, 10431, 11414, 9499, 9880, 9050, 4065, 4630, 3863, 944, 0, 68, 0, 17, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 54, 0, 177, 0, 1496, 3565, 2765, 7482, 9672, 8491, 9962, 9239, 8673, 8831, 8836, 7985, 8552, 9862, 9951, 10391, 10050, 10047, 10554, 9052, 11376, 5072, 0, 630, 0, 181, 0, 36, 0, 0, 0, 0, 0, 0, 4, 0, 19, 0, 77, 0, 730, 2077, 2334, 2196, 5261, 7076, 6654, 6856, 7252, 2916, 0, 346, 0, 97, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 1, 1, 0, 1, 236, 1936, 980, 0, 0, 959, 2092, 4655, 7907, 8302, 8741, 8651, 9472, 9059, 9076, 3312, 0, 377, 0, 108, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 21, 0, 89, 0, 859, 2726, 3752, 3184, 5818, 9019, 7876, 8559, 7863, 8501, 3583, 0, 390, 0, 0, 301, 0, 2907, 6319, 6001, 6089, 7270, 3472, 0, 442, 0, 123, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 74, 0, 259, 0, 2200, 5623, 5588, 6342, 6507, 6843, 7331, 7920, 8261, 8792, 9129, 9177, 9382, 9362, 9430, 9868, 8925, 8426, 8163, 7743, 8483, 4665, 363, 30, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 15, 0, 49, 0, 439, 967, 248, 18, 748, 954, 3118, 5568, 6359, 6702, 6398, 6548, 2308, 0, 222, 0, 65, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 13, 0, 44, 0, 391, 951, 269, 0, 22, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 57, 0, 215, 0, 1691, 3437, 2728, 1905, 4455, 7603, 7206, 6101, 2428, 588, 143, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 52, 0, 191, 0, 1717, 3745, 3513, 1485, 0, 186, 0, 46, 0, 0, 12, 0, 59, 0, 909, 3985, 4054, 2704, 7296, 13354, 16307, 16995, 17131, 17726, 17787, 18257, 17705, 18155, 16963, 17209, 15931, 8220, 9602, 11344, 8179, 8209, 8445, 8820, 8448, 7912, 5082, 2060, 2505, 3541, 3275, 2969, 3239, 2862, 2562, 2602, 2669, 2471, 2932, 1322, 0, 1345, 7455, 5619, 0, 258, 0, 89, 0, 55, 0, 145, 0, 1531, 5428, 7453, 8431, 9042, 5685, 3893, 8038, 9815, 9982, 9170, 5810, 1327, 0, 111, 0, 30, 0, 7, 0, 2, 0, 130, 841, 1007, 748, 910, 712, 1020, 459, 2034, 1928, 0, 1749, 1483, 771, 1313, 2083, 1018, 0, 129, 0, 33, 0, 0, 26, 0, 99, 0, 811, 1698, 363, 0, 8, 7, 0, 211, 794, 751, 305, 142, 264, 109, 0, 12, 0, 3, 0, 14, 0, 64, 0, 241, 0, 2465, 8492, 11189, 9774, 11571, 8205, 2394, 1328, 0, 190, 0, 0, 866, 5164, 7119, 5653, 7604, 9420, 9764, 8637, 6121, 1945, 0, 210, 0, 53, 0, 0, 63, 0, 251, 0, 1650, 1650, 0, 251, 0, 68, 0, 0, 37, 0, 144, 0, 997, 1244, 0, 1130, 1941, 1876, 613, 0, 0, 116, 0, 1357, 3654, 3092, 3638, 3566, 3885, 3406, 3487, 1723, 0, 354, 0, 1111, 2379, 2996, 2161, 617, 666, 53, 11, 0, 0, 0, 0, 0, 0, 0, 49, 0, 244, 0, 863, 0, 6982, 16187, 13908, 16086, 17402, 17858, 8401, 0, 4496, 11285, 12036, 12616, 12593, 13259, 13274, 13410, 12962, 14533, 14271, 13558, 11948, 9084, 3223, 0, 313, 0, 0, 869, 2961, 2531, 3780, 863, 1603, 2154, 0, 354, 0, 84, 0, 0, 44, 0, 194, 0, 2532, 11965, 18646, 12237, 7713, 11216, 10278, 11879, 14209, 14469, 14582, 13890, 14304, 7517, 385, 78, 0, 0, 583, 614, 0, 88, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 33, 0, 114, 0, 1572, 7010, 9175, 10119, 13892, 15871, 15533, 15244, 15244, 15068, 15186, 15672, 15960, 16090, 16159, 16240, 16264, 16261, 16882, 16523, 17268, 14255, 10708, 6180, 0, 1284, 1012, 0, 144, 0, 44, 0, 9, 0, 0, 0, 0, 0, 71, 0, 349, 0, 1215, 0, 9947, 23315, 19759, 22169, 21483, 22462, 23550, 22784, 23442, 20618, 19133, 18552, 19496, 13813, 5780, 6143, 6946, 10433, 5076, 2389, 6158, 7825, 6253, 7414, 10198, 8479, 8814, 8012, 7002, 8817, 11815, 8771, 5517, 7638, 8760, 9562, 11922, 13938, 14100, 14057, 14199, 13885, 14492, 13328, 16218, 12856, 7435, 9603, 7932, 7983, 8664, 9986, 8482, 12333, 11731, 10081, 15530, 15897, 16584, 16863, 17089, 17005, 16572, 15465, 15806, 14840, 15957, 8129, 2403, 2322, 0, 391, 0, 97, 0, 12, 0, 0, 0, 0, 0, 0, 43, 0, 217, 0, 772, 0, 6266, 14342, 12805, 11127, 9810, 4278, 0, 1263, 0, 241, 0, 23, 41, 0, 255, 0, 2208, 6066, 7001, 2814, 0, 336, 0, 94, 0, 10, 7, 0, 90, 0, 329, 0, 2705, 6841, 8859, 11125, 11726, 12121, 11304, 11737, 11281, 11951, 10799, 13046, 5744, 0, 619, 225, 3837, 6336, 6342, 5480, 6503, 8303, 8939, 8834, 8936, 8994, 10528, 9334, 3353, 113, 43, 0, 18, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 87, 0, 305, 0, 2463, 5520, 4688, 4900, 5180, 4288, 6194, 1142, 3719, 4827, 0, 1103, 0, 3381, 8276, 2683, 0, 247, 0, 81, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 22, 0, 64, 0, 577, 1094, 0, 2982, 7408, 7091, 7293, 7088, 7181, 7149, 7132, 7201, 7048, 7448, 7629, 9344, 10193, 11681, 13605, 13155, 12041, 10455, 4077, 0, 684, 0, 104, 0, 21, 0, 0, 0, 0, 2, 0, 33, 0, 152, 130, 3003, 4813, 7427, 10188, 10373, 10647, 13119, 14856, 17002, 11536, 2706, 1980, 1116, 1498, 1282, 1432, 1270, 1541, 682, 0, 84, 0, 29, 0, 27, 0, 77, 0, 2009, 9429, 13803, 15597, 18894, 20121, 18468, 18383, 13849, 12849, 13886, 11045, 12398, 10085, 9213, 10950, 11292, 13389, 14416, 13192, 15303, 12920, 8698, 10266, 13933, 15641, 9507, 5910, 6671, 6241, 6533, 6281, 6583, 6057, 7951, 11585, 12634, 13873, 14663, 15053, 15023, 16230, 16152, 13907, 5224, 0, 391, 0, 106, 0, 8, 4, 0, 463, 2268, 1404, 1167, 3889, 3452, 5350, 9478, 12845, 14243, 14695, 13193, 11740, 10385, 11662, 14723, 14773, 15928, 16158, 16284, 16410, 16043, 16772, 15412, 18172, 8565, 0, 4931, 9861, 4731, 3987, 8831, 8898, 10891, 4283, 0, 515, 0, 2310, 5965, 3314, 4240, 8324, 8031, 7625, 6684, 6353, 4052, 4637, 7923, 8768, 9096, 10078, 10896, 12887, 15706, 17267, 17282, 11844, 7764, 4894, 3652, 5652, 5124, 5572, 5096, 5782, 4525, 8585, 12917, 12682, 14371, 13360, 12917, 11590, 11113, 4830, 0, 349, 0, 103, 0, 29, 0, 49, 0, 292, 114, 326, 1273, 4055, 5732, 1804, 794, 2713, 3124, 2338, 691, 0, 1196, 4477, 9250, 4039, 0, 2099, 2944, 6662, 7883, 7457, 7964, 7155, 8675, 3815, 0, 439, 0, 10, 153, 0, 2125, 7270, 11311, 13367, 12986, 13651, 13223, 14025, 14171, 13848, 12538, 12206, 12055, 10446, 11739, 12602, 12990, 13182, 12851, 11080, 13799, 6067, 0, 866, 0, 1425, 3721, 4190, 4798, 5137, 5585, 6753, 7034, 7000, 6991, 7035, 6968, 6600, 2192, 0, 235, 0, 68, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3563, 4912, 3282, 6004, 0, 16308, 35204, 28494, 32052, 30323, 31440, 31312, 31580, 31495, 31532, 31477, 31585, 31370, 32071, 32792, 32304, 31661, 30746, 25671, 14537, 14863, 21251, 22270, 23832, 23247, 23420, 23942, 23873, 24316, 24608, 24231, 24216, 23556, 22911, 22693, 21145, 21162, 21477, 21751, 21454, 21694, 21995, 23006, 22307, 22824, 8504, 0, 1458, 0, 357, 0, 78, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 168, 0, 554, 0, 4753, 11012, 2899, 0, 220, 0, 78, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 100, 0, 334, 0, 2931, 7863, 6507, 6245, 3618, 1199, 1853, 1333, 1318, 947, 2876, 2054, 4814, 11458, 13159, 11160, 8622, 6763, 6117, 9283, 10269, 11479, 11506, 10540, 10626, 9999, 10601, 10991, 10659, 5862, 1030, 853, 1887, 6671, 3221, 0, 400, 0, 165, 0, 250, 0, 779, 0, 6076, 12502, 8390, 9673, 8993, 9456, 9221, 9492, 10683, 10357, 10102, 10775, 10179, 9873, 9161, 8621, 9109, 9318, 9936, 10152, 10426, 10838, 11005, 10674, 9365, 7198, 3142, 1570, 646, 265, 967, 4551, 7843, 8911, 8063, 6816, 8208, 7811, 9050, 9566, 9481, 9461, 9584, 9285, 10201, 10299, 9629, 9611, 9227, 9576, 9516, 9810, 9057, 8558, 7876, 7186, 7311, 7445, 7454, 7121, 7407, 7607, 7610, 7656, 7662, 7726, 7552, 7390, 7537, 8002, 7240, 7129, 7372, 8501, 3510, 0, 421, 0, 120, 0, 24, 0, 48, 0, 240, 0, 842, 0, 6765, 15236, 12775, 13773, 12837, 13326, 13399, 13406, 13220, 14061, 13343, 13789, 11671, 11178, 4780, 0, 594, 0, 166, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 212, 0, 746, 0, 6000, 13500, 11389, 12800, 13024, 13806, 13320, 13414, 11764, 10477, 10457, 9969, 10122, 9589, 8989, 9471, 10141, 9969, 9748, 9371, 10258, 3996, 0, 493, 0, 230, 0, 701, 916, 0, 67, 0, 17, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 77, 0, 276, 0, 1803, 1829, 0, 393, 0, 445, 0, 8245, 13430, 9614, 11104, 8475, 7399, 9377, 8406, 8793, 3413, 0, 404, 0, 119, 0, 33, 0, 35, 0, 309, 915, 1194, 1349, 1586, 2240, 1525, 450, 424, 2102, 5449, 6586, 6405, 6354, 6618, 6039, 7254, 3216, 0, 399, 0, 114, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 60, 0, 213, 0, 1761, 5113, 8189, 11435, 7619, 7764, 10205, 9527, 9881, 9638, 9738, 9728, 9661, 9813, 9523, 10228, 8251, 1842, 0, 135, 0, 41, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 75, 0, 263, 0, 2109, 4817, 3920, 4490, 3978, 4607, 3528, 7209, 11237, 3228, 0, 0, 1369, 5541, 7074, 8967, 9885, 11353, 7656, 3477, 3091, 2823, 2354, 2100, 3525, 4217, 2644, 204, 21, 0, 8, 0, 1, 0, 8, 0, 38, 0, 412, 1647, 2935, 4398, 5024, 6794, 9502, 10195, 10058, 10142, 10053, 10178, 9950, 10728, 11822, 11383, 11235, 10637, 9831, 9785, 9719, 10095, 9703, 9485, 10245, 9262, 4470, 2750, 1485, 0, 208, 0, 56, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 53, 0, 191, 0, 1587, 3999, 4466, 5233, 5135, 5521, 5731, 6096, 7043, 7551, 7425, 7464, 7482, 7401, 7588, 6975, 6491, 6672, 6554, 7105, 6499, 6177, 7148, 7141, 7298, 6989, 3913, 660, 0, 35, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 23, 0, 74, 0, 739, 2140, 747, 0, 75, 0, 24, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 24, 0, 87, 0, 727, 1807, 1792, 2160, 2173, 2205, 2162, 2231, 2107, 2359, 1456, 78, 25, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 24, 0, 63, 0, 546, 1552, 2253, 3333, 4022, 4770, 5867, 6163, 6142, 5885, 5827, 6281, 6473, 6478, 5863, 5642, 5753, 5581, 5886, 5333, 6430, 2843, 0, 353, 0, 101, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 53, 0, 223, 0, 1343, 1455, 4607, 4345, 1366, 967, 649, 2368, 1403, 1848, 1604, 1758, 1620, 1823, 1200, 470, 460, 15, 209, 825, 750, 364, 333, 479, 196, 0, 23, 0, 6, 0, 3, 0, 7, 0, 110, 467, 836, 1100, 1473, 966, 2533, 4244, 4630, 5689, 6550, 6113, 6005, 6175, 5748, 6731, 6803, 6280, 6083, 6190, 6015, 6337, 5745, 6924, 3062, 0, 380, 0, 108, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 60, 0, 220, 0, 1455, 1826, 1885, 4520, 4701, 5045, 5056, 4566, 3593, 3708, 2190, 162, 20, 0, 8, 0, 0, 4, 0, 11, 0, 212, 864, 396, 0, 47, 0, 14, 0, 3, 0, 1, 0, 0, 1, 0, 0, 542, 4523, 6811, 6684, 8056, 6459, 6650, 7038, 6724, 8393, 7793, 7398, 8325, 7639, 7453, 7493, 7264, 6936, 5452, 5315, 4931, 4513, 4695, 4508, 4778, 4326, 5201, 2351, 0, 272, 0, 78, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 83, 0, 316, 0, 2826, 3451, 4772, 6054, 3688, 5184, 6522, 5310, 4918, 2048, 84, 97, 2154, 5656, 4550, 5001, 4951, 4633, 5504, 2451, 0, 303, 0, 84, 0, 7, 4, 0, 46, 0, 541, 2412, 4736, 7388, 8458, 8399, 8865, 9308, 8894, 8634, 8122, 6963, 6750, 7345, 8718, 8414, 7501, 7620, 7985, 8293, 7977, 7105, 7453, 7353, 7951, 6337, 3670, 4003, 3801, 3835, 3965, 3625, 4355, 1927, 0, 239, 0, 68, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 10, 0, 154, 407, 26, 2688, 6221, 6270, 7136, 2827, 0, 336, 0, 99, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 11, 0, 45, 0, 1040, 6450, 11058, 12277, 13058, 12929, 11676, 12297, 9750, 7685, 7992, 5196, 1413, 0, 135, 0, 34, 0, 6, 0, 0, 0, 0, 0, 0, 14, 0, 76, 0, 277, 0, 2124, 4501, 5299, 7614, 7499, 7223, 7919, 9213, 9772, 8852, 6956, 6721, 5955, 5781, 6941, 6361, 7545, 8839, 8581, 8763, 8736, 8718, 8222, 8730, 7736, 8136, 3331, 0, 402, 0, 115, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 31, 0, 204, 204, 0, 31, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 45, 0, 156, 0, 1620, 5586, 6717, 7843, 9627, 9007, 8443, 7346, 5764, 5068, 3953, 4964, 6181, 6213, 6205, 6315, 6387, 6841, 7680, 8569, 9153, 8476, 7717, 8860, 9585, 8093, 7871, 3706, 0, 206, 0, 45, 0, 0, 116, 0, 938, 1600, 240, 0, 139, 0, 1342, 4050, 5539, 7065, 7498, 8177, 9187, 9908, 9877, 10050, 9732, 9461, 8985, 8919, 7949, 8086, 7602, 8548, 3914, 0, 601, 0, 525, 0, 3114, 6920, 6018, 6375, 5561, 6145, 5313, 4026, 3760, 3846, 3715, 3952, 3468, 5226, 8071, 8224, 8484, 9377, 9353, 10005, 10925, 11375, 13425, 9593, 5668, 6603, 5843, 6238, 6503, 6222, 6492, 6745, 6662, 7448, 7885, 7917, 9220, 10207, 9676, 9311, 9810, 8938, 9554, 6118, 705, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 252, 2760, 7381, 8972, 10749, 12075, 12189, 12913, 13168, 11229, 8852, 10085, 9913, 11392, 4556, 0, 394, 0, 0, 2236, 5550, 6860, 3221, 0, 564, 0, 69, 0, 0, 113, 116, 0, 17, 0, 23, 0, 103, 0, 378, 0, 2982, 7312, 10758, 15637, 15309, 15307, 13428, 12876, 13746, 12231, 8612, 6452, 6488, 6540, 6636, 8169, 9144, 9151, 9081, 9363, 10272, 11248, 12059, 13071, 12939, 12025, 11273, 6897, 1468, 0, 110, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 10, 0, 86, 0, 352, 0, 1808, 6, 4508, 12793, 12762, 14554, 14153, 15185, 15164, 14704, 14781, 13539, 12217, 13563, 9237, 2841, 2500, 893, 0, 95, 0, 30, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 230, 0, 804, 0, 6489, 14758, 12315, 13399, 12580, 12960, 12531, 8313, 5848, 6235, 6552, 5809, 9033, 12112, 10474, 10691, 10273, 10849, 9928, 10748, 11440, 10181, 10126, 10638, 10225, 3110, 0, 313, 0, 92, 0, 20, 0, 0, 0, 0, 0, 0, 53, 0, 264, 0, 924, 0, 7405, 16609, 13758, 15362, 14026, 14980, 14821, 14434, 11630, 9496, 10199, 10608, 10018, 8782, 8769, 8604, 8455, 8549, 8233, 7319, 8170, 8107, 8947, 4297, 0, 1118, 1173, 6921, 6249, 4088, 3341, 0, 6006, 8853, 10403, 9991, 9134, 11452, 11099, 11371, 11208, 11332, 11175, 11457, 10708, 10933, 10759, 11552, 7964, 5249, 5972, 7715, 11179, 10109, 10350, 10351, 10226, 10646, 10510, 11027, 9783, 9462, 6422, 5852, 3205, 0, 441, 0, 120, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 158, 0, 552, 0, 4326, 9218, 7465, 8511, 5873, 1583, 0, 145, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 41, 0, 336, 961, 1871, 2512, 2268, 2495, 2177, 2703, 1717, 4566, 4967, 1777, 2598, 1739, 3058, 4730, 4260, 3052, 3075, 3228, 3333, 1375, 0, 166, 0, 46, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8841, 8746, 8917, 8357, 8333, 8129, 9581, 6788, 10260, 0, 18539, 25962, 8270, 10188, 6543, 10222, 10324, 5212, 0, 430, 75, 0, 3599, 9304, 8538, 9130, 8907, 8986, 8788, 8728, 8559, 7809, 7477, 7500, 7953, 8656, 8754, 8960, 9167, 9412, 9476, 9475, 9446, 9531, 9348, 9715, 8957, 11306, 13197, 12987, 4931, 0, 599, 0, 280, 0, 453, 0, 3311, 7424, 7622, 8885, 8255, 10473, 11369, 11620, 12415, 12016, 11591, 11677, 12052, 12274, 12311, 12221, 12061, 12328, 12342, 11268, 10102, 11120, 9505, 8422, 8667, 8745, 8883, 8044, 8432, 8091, 8535, 7815, 9200, 4693, 178, 1819, 1297, 1469, 1237, 1606, 1940, 2228, 2780, 3005, 3000, 2850, 2677, 2650, 2752, 2706, 2931, 2145, 1108, 1328, 2244, 3185, 2690, 3207, 2173, 160, 27, 0, 26, 0, 56, 0, 1102, 1777, 1843, 2568, 1935, 1580, 1646, 1650, 1582, 1743, 1396, 2582, 3960, 3802, 4046, 4054, 4208, 4265, 4304, 4327, 4482, 4068, 3962, 4270, 4182, 4231, 4209, 4234, 4336, 4411, 4430, 4441, 4435, 4458, 4463, 4398, 4410, 4399, 4422, 4503, 4540, 4448, 4388, 4408, 4396, 4202, 3994, 3766, 3543, 3537, 3535, 3533, 3536, 3538, 3531, 3430, 2863, 3741, 1672, 0, 207, 0, 59, 0, 12, 0, 3, 0, 12, 0, 37, 0, 524, 2317, 2678, 3327, 4198, 4087, 4106, 3967, 3713, 3766, 3713, 3528, 4020, 3819, 3731, 3541, 3905, 1606, 0, 193, 0, 55, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 35, 0, 122, 0, 1130, 3337, 3484, 3532, 3625, 3536, 3523, 944, 499, 1984, 2771, 1442, 0, 189, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 36, 0, 121, 0, 1014, 2240, 542, 0, 36, 0, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 149, 0, 527, 0, 3994, 7752, 5631, 6344, 5306, 6697, 7001, 6842, 7333, 6593, 6097, 5256, 3991, 4157, 3122, 2320, 1317, 196, 358, 113, 0, 10, 0, 2, 0, 4, 0, 24, 0, 136, 518, 2941, 4074, 2630, 1692, 358, 0, 28, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 37, 0, 337, 1243, 2889, 3822, 3508, 3767, 3436, 3970, 2959, 6051, 8009, 6849, 7351, 6492, 4059, 3596, 4879, 4712, 4998, 5713, 4051, 3799, 2155, 0, 299, 0, 82, 0, 14, 0, 0, 0, 0, 0, 1, 0, 4, 0, 164, 1333, 2785, 3363, 2589, 3645, 4544, 5340, 6551, 6388, 6363, 6616, 6037, 7255, 3213, 0, 399, 0, 114, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 47, 0, 175, 0, 1267, 2324, 2553, 2159, 677, 1375, 713, 1618, 5, 5117, 10251, 8376, 8137, 2344, 0, 231, 0, 75, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 43, 0, 148, 0, 1417, 4353, 4737, 4631, 4852, 4410, 5312, 2349, 0, 290, 0, 74, 0, 0, 65, 0, 530, 1004, 1110, 599, 0, 81, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 315, 1581, 3441, 4812, 6261, 7046, 6820, 6946, 6850, 6953, 6794, 7221, 7270, 6755, 6287, 5468, 4667, 4875, 4802, 4630, 7006, 2899, 0, 342, 0, 101, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 16, 0, 57, 0, 1426, 1857, 1841, 3189, 3595, 2206, 224, 17, 62, 1366, 2219, 2000, 2066, 2106, 1944, 2323, 1032, 0, 127, 0, 36, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 35, 0, 122, 0, 1341, 5183, 7102, 6852, 5963, 6631, 8708, 9171, 8230, 7598, 7434, 6949, 6400, 6645, 6388, 6768, 6119, 7384, 3265, 0, 405, 0, 116, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 85, 0, 304, 0, 2537, 6626, 7970, 8345, 6176, 4938, 4580, 5743, 7663, 8038, 7498, 6716, 7750, 3333, 0, 408, 0, 116, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 158, 0, 551, 0, 4578, 10872, 7699, 2688, 0, 256, 0, 52, 0, 0, 84, 0, 775, 2202, 3620, 4268, 3485, 3181, 3730, 5238, 7707, 8467, 7843, 8025, 8035, 7837, 8300, 7319, 10549, 13472, 12174, 13140, 14252, 14030, 13693, 14032, 13728, 13491, 14188, 11319, 9089, 9451, 7779, 7692, 6721, 5517, 5232, 6374, 6766, 6615, 6552, 5623, 4746, 4312, 3305, 4013, 1930, 0, 247, 0, 70, 0, 14, 0, 0, 0, 6, 0, 28, 0, 83, 0, 981, 4016, 4412, 5016, 2156, 0, 268, 0, 77, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 35, 0, 278, 1136, 3592, 1873, 0, 241, 0, 65, 0, 0, 49, 0, 197, 0, 1601, 3807, 3920, 4551, 4353, 4364, 4527, 4133, 4967, 2199, 0, 273, 0, 78, 0, 14, 0, 0, 0, 3, 0, 2, 206, 2152, 3659, 3419, 2486, 2299, 3518, 4035, 4204, 4014, 1285, 0, 133, 0, 39, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 30, 0, 99, 0, 1798, 9704, 13268, 12855, 13134, 13442, 11422, 8819, 6551, 4087, 4449, 3772, 4275, 4280, 6268, 8852, 8781, 8799, 8582, 8400, 9809, 10349, 3004, 0, 0, 1531, 5581, 6772, 7458, 7602, 7780, 7813, 7633, 8021, 7281, 8768, 3880, 0, 527, 0, 349, 0, 750, 0, 5754, 12038, 5598, 4378, 3333, 3101, 2431, 2896, 1759, 364, 332, 1853, 3881, 4179, 3463, 6521, 8218, 5493, 10531, 4865, 0, 765, 2917, 7730, 8979, 9197, 10286, 9121, 10435, 7736, 3783, 4951, 4535, 4442, 5148, 2327, 0, 286, 0, 81, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 7, 155, 2353, 6624, 9378, 11832, 11006, 8787, 8485, 8160, 8580, 8420, 8538, 8716, 8674, 8711, 8671, 8733, 8620, 8921, 8925, 8464, 5330, 868, 0, 36, 0, 11, 0, 19, 0, 39, 0, 62, 0, 1805, 9129, 2762, 3336, 10134, 7031, 7210, 8841, 11611, 12251, 12547, 12767, 11623, 11479, 12965, 13796, 13274, 15523, 8814, 6659, 14528, 6535, 100, 129, 0, 0, 147, 0, 1613, 4457, 7932, 9379, 9933, 6722, 3703, 7798, 3843, 5017, 8629, 8598, 8661, 6920, 7280, 7400, 7548, 7598, 7781, 7397, 7832, 8337, 8566, 8982, 10387, 9754, 7897, 8021, 7844, 8264, 6521, 5141, 6498, 7650, 8169, 8016, 8143, 8266, 8306, 8332, 8330, 8320, 8345, 8297, 8421, 8266, 7622, 7610, 7230, 7042, 4056, 1517, 2374, 2624, 2811, 2722, 2005, 558, 443, 543, 64, 23, 0, 0, 34, 0, 123, 0, 1170, 2971, 2580, 3589, 3746, 776, 2033, 1688, 0, 252, 0, 71, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 50, 160, 2480, 2452, 2741, 5826, 5899, 6283, 6860, 7436, 7214, 6416, 5828, 7519, 3210, 0, 205, 134, 0, 2896, 7387, 7011, 7239, 6860, 7290, 6943, 6772, 6891, 6687, 7051, 6389, 7703, 3407, 0, 423, 0, 121, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 35, 0, 125, 0, 819, 819, 0, 125, 0, 35, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 32, 0, 97, 0, 1353, 5682, 4577, 2676, 3642, 3920, 3871, 3459, 4249, 4171, 4294, 5915, 5358, 4516, 3665, 838, 0, 62, 0, 17, 0, 0, 14, 0, 66, 0, 593, 2071, 3214, 4844, 4465, 5067, 2352, 0, 3519, 2165, 5107, 8845, 10038, 4557, 0, 579, 0, 160, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 211, 0, 734, 0, 5908, 13182, 10064, 10949, 10361, 10566, 10213, 10247, 9775, 9074, 3144, 0, 347, 0, 86, 399, 3750, 4842, 5317, 5142, 3906, 4590, 4419, 4430, 5179, 4844, 5378, 6588, 6348, 6911, 6914, 7054, 6617, 6383, 5136, 1222, 0, 98, 0, 29, 0, 15, 0, 44, 0, 154, 0, 1016, 1052, 0, 228, 0, 752, 2055, 1425, 2686, 4408, 4498, 5662, 7318, 8062, 8484, 9396, 9763, 9897, 10390, 9665, 9674, 9206, 6973, 2091, 0, 69, 341, 381, 31, 0, 1398, 3758, 1191, 0, 112, 0, 37, 0, 5, 3, 0, 46, 0, 161, 0, 2176, 5036, 5460, 5943, 6313, 7355, 8191, 9081, 8949, 7696, 6751, 7102, 3852, 2907, 4410, 3943, 4438, 4088, 4230, 5967, 7015, 6242, 6113, 6163, 6052, 6298, 5441, 5308, 2087, 0, 248, 0, 70, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 160, 0, 560, 0, 4753, 12149, 11734, 12559, 12102, 12346, 12197, 12325, 12153, 12481, 11376, 10126, 9872, 9514, 8271, 7743, 2963, 0, 329, 0, 31, 67, 0, 896, 1709, 1410, 2091, 2095, 2866, 3388, 3654, 3929, 3545, 3894, 3175, 3183, 1479, 0, 190, 0, 53, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21409, 19859, 22667, 13535, 3355, 6731, 5552, 7025, 4020, 344, 354, 0, 52, 0, 0, 111, 82, 4584, 9199, 8580, 12465, 15412, 15115, 13887, 19365, 22735, 21621, 21980, 23198, 26349, 35888, 15774, 0, 1766, 1844, 0, 15676, 35875, 28870, 31443, 29537, 29685, 29213, 29354, 29334, 29295, 29385, 28802, 27180, 30073, 33573, 30196, 26211, 24561, 27386, 30100, 29864, 30357, 31334, 31248, 31249, 29373, 27577, 26913, 26677, 24346, 20622, 18135, 22780, 27090, 25969, 25514, 18210, 6850, 2596, 3745, 2840, 2725, 3624, 4372, 3611, 2616, 3092, 3443, 2945, 3125, 3064, 3034, 3166, 2883, 3469, 1535, 0, 190, 0, 54, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 222, 1972, 4177, 3871, 1716, 9971, 17813, 19890, 22497, 25263, 29247, 30765, 31766, 32014, 32570, 32606, 32543, 32410, 30411, 29553, 27197, 24051, 19653, 20244, 11871, 2700, 8062, 13570, 12267, 6861, 6696, 4904, 2115, 1185, 1675, 1656, 1878, 1790, 1841, 1809, 1837, 1800, 1900, 1929, 1819, 1798, 1644, 2000, 2058, 1504, 1628, 1207, 298, 0, 478, 1296, 1920, 2736, 2793, 2879, 2756, 2421, 2189, 3874, 11592, 16299, 16613, 17135, 17693, 7777, 0, 2804, 4905, 4572, 6537, 4349, 0, 242, 0, 75, 0, 11, 0, 0, 0, 0, 0, 20, 0, 96, 0, 355, 0, 3276, 9408, 10650, 9941, 14931, 17336, 17111, 19869, 19464, 20097, 20030, 21149, 21372, 21300, 21140, 20917, 20892, 20472, 21495, 21777, 21193, 20451, 20070, 20388, 19645, 19269, 18944, 19056, 19541, 20121, 21614, 22239, 22230, 21966, 22582, 21386, 23803, 15686, 6590, 9275, 5820, 5898, 4986, 10205, 15356, 14837, 17379, 14549, 12999, 18290, 7522, 0, 883, 0, 258, 0, 45, 0, 0, 79, 0, 518, 520, 0, 88, 0, 42, 46, 1191, 2081, 638, 0, 59, 0, 19, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 2, 0, 56, 0, 177, 390, 6797, 4338, 0, 680, 0, 593, 0, 1493, 0, 11697, 26562, 20746, 20119, 12511, 11461, 7436, 2720, 4886, 4745, 4968, 3231, 1875, 2305, 1512, 383, 0, 32, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 17, 0, 79, 0, 1038, 5017, 8937, 3372, 0, 0, 1439, 2161, 0, 203, 0, 50, 0, 8, 0, 0, 0, 44, 0, 231, 0, 819, 0, 6701, 16371, 18164, 24837, 25997, 26852, 27183, 27058, 27071, 27171, 26891, 27456, 26320, 29711, 30861, 28563, 29622, 28824, 28270, 26928, 26788, 25090, 23674, 21282, 19242, 19662, 18696, 18251, 17643, 17359, 19582, 23296, 29065, 24491, 18128, 20036, 20324, 20072, 18404, 18582, 16621, 17329, 20745, 21985, 23786, 26980, 30248, 27207, 24655, 8621, 0, 967, 0, 278, 0, 56, 0, 0, 8, 0, 50, 0, 184, 0, 1370, 3044, 3986, 5719, 3721, 4408, 2166, 0, 286, 0, 82, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 0, 74, 0, 529, 606, 0, 219, 0, 2397, 12691, 17874, 18698, 19780, 21679, 23784, 25551, 28376, 28516, 29088, 27641, 25858, 18182, 13675, 7840, 2615, 2044, 0, 2316, 2542, 2636, 2542, 2677, 2440, 2930, 1300, 0, 161, 0, 46, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 115, 0, 426, 0, 3324, 7323, 7771, 6469, 5401, 9081, 8198, 15687, 13748, 7461, 9655, 8347, 9386, 8232, 10078, 4427, 0, 551, 0, 157, 0, 32, 0, 0, 41, 0, 211, 0, 633, 0, 6143, 20858, 23005, 35752, 16749, 0, 2170, 155, 0, 1864, 0, 16200, 35887, 28411, 28820, 24897, 25807, 25584, 24682, 23394, 22962, 21977, 21060, 20947, 20918, 20986, 20870, 21066, 20662, 22491, 26918, 24938, 24512, 26294, 27118, 28057, 26810, 26861, 25879, 25380, 25728, 25930, 24681, 25147, 22961, 26533, 29279, 28322, 20773, 15121, 17157, 15156, 5694, 0, 754, 0, 324, 178, 102, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 1, 5, 0, 65, 250, 3571, 1263, 571, 0, 8862, 22708, 22940, 26001, 26565, 28984, 29765, 30587, 30369, 30229, 28155, 27027, 21821, 20957, 10807, 1577, 6606, 11552, 13592, 17006, 8168, 0, 1544, 2036, 5143, 5295, 4866, 4985, 5852, 4827, 4042, 4630, 4166, 4038, 4231, 4090, 4286, 3960, 4585, 2579, 563, 654, 0, 69, 0, 22, 0, 34, 0, 117, 0, 987, 2458, 2175, 2725, 2745, 2649, 1892, 1761, 5779, 16148, 6200, 1397, 4069, 0, 1546, 3764, 2274, 0, 287, 0, 77, 0, 17, 0, 0, 0, 0, 31, 0, 152, 0, 399, 0, 4135, 15416, 13907, 32491, 15305, 0, 0, 21626, 16844, 9885, 40071, 28345, 32989, 26419, 25433, 24643, 23160, 23512, 23164, 22261, 21730, 20848, 19990, 17846, 17124, 16946, 17101, 16723, 15832, 15303, 14681, 13335, 17082, 19091, 18862, 11418, 5711, 7839, 6869, 7346, 7154, 7156, 7333, 6635, 7015, 10690, 8157, 10144, 15435, 6961, 1885, 3353, 1344, 47, 9, 0, 9, 0, 3, 0, 0, 0, 4, 0, 46, 0, 176, 0, 2708, 3195, 4164, 3050, 0, 309, 0, 85, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 2, 0, 114, 1030, 2547, 1013, 0, 0, 259, 0, 3786, 15076, 19188, 20456, 24418, 30628, 33129, 32643, 32603, 33112, 31922, 34441, 26054, 15280, 7960, 1968, 9038, 10337, 13979, 6522, 0, 766, 0, 223, 0, 44, 0, 0, 0, 0, 0, 3, 0, 18, 0, 66, 0, 647, 2168, 2833, 2846, 2349, 755, 0, 80, 0, 23, 0, 4, 0, 11, 0, 49, 0, 161, 0, 1753, 6618, 6309, 6330, 6061, 10020, 5943, 0, 613, 0, 373, 124, 0, 19, 0, 8, 0, 1, 0, 0, 0, 0, 0, 3, 0, 41, 0, 1050, 8371, 21608, 28772, 25799, 24174, 24978, 27127, 29390, 29552, 29548, 29342, 29435, 29356, 29468, 29277, 29657, 28352, 26349, 24994, 23775, 21184, 16997, 15475, 16514, 17047, 20513, 22581, 21707, 21185, 20123, 18854, 19355, 13636, 9362, 10885, 11465, 11738, 10515, 11621, 11095, 11364, 11047, 11000, 6352, 4774, 19842, 27324, 24961, 22807, 19838, 15647, 16925, 7889, 0, 2028, 547, 1320, 957, 1059, 1172, 552, 0, 129, 0, 430, 401, 0, 61, 0, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 32, 0, 111, 0, 953, 2551, 2428, 1954, 475, 0, 30, 0, 0, 60, 0, 188, 0, 2543, 9750, 4259, 0, 559, 0, 545, 474, 0, 708, 1777, 8661, 5080, 0, 683, 0, 198, 0, 40, 0, 2, 0, 11, 0, 33, 0, 788, 2022, 1930, 2340, 2803, 2092, 1026, 629, 274, 0, 14, 18, 0, 151, 0, 1229, 2496, 2878, 1857, 5799, 10307, 9362, 9969, 7102, 5630, 5062, 4607, 5049, 5320, 4426, 2888, 3594, 2016, 902, 1473, 1242, 1385, 1281, 1384, 1242, 1498, 646, 0, 0, 191, 0, 925, 0, 11595, 20859, 31334, 17556, 0, 4993, 1337, 3698, 1047, 4066, 0, 14244, 31776, 26070, 28522, 26770, 27015, 26476, 26684, 26459, 26093, 25929, 26107, 26100, 25807, 25852, 25993, 26227, 25976, 26774, 26882, 26198, 26382, 26399, 26187, 26674, 25643, 29110, 32806, 31548, 31826, 31462, 31948, 31570, 32330, 30749, 27840, 27005, 23391, 20387, 16294, 4800, 0, 1053, 702, 1450, 1988, 1581, 1948, 807, 1616, 2808, 1263, 2841, 2799, 2130, 937, 0, 367, 8, 18, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 62, 0, 219, 0, 1737, 3791, 3182, 3796, 3760, 3595, 4133, 2961, 5220, 913, 12028, 7018, 5640, 27766, 23454, 34095, 16727, 0, 5156, 0, 15335, 30414, 22549, 24093, 19979, 22695, 19527, 15421, 17872, 18051, 17987, 17647, 14236, 16172, 8600, 4278, 5379, 1348, 3175, 2624, 3427, 3196, 2275, 1878, 1617, 1391, 1444, 1431, 1571, 1274, 1881, 725, 2869, 0, 12716, 27405, 24017, 26393, 26632, 28518, 28593, 29176, 29517, 29398, 27785, 29535, 30825, 32743, 30294, 36382, 17423, 0, 4912, 0, 16386, 36837, 26364, 33879, 12795, 0, 4282, 0, 904, 0, 209, 0, 0, 46, 0, 185, 0, 1590, 3135, 3272, 2200, 4566, 0, 16189, 33521, 29194, 32075, 30224, 30953, 30040, 29855, 26267, 25580, 30358, 29411, 24873, 22835, 22887, 22385, 21956, 21924, 21027, 21571, 18309, 16807, 10285, 3842, 6330, 6278, 6699, 5699, 5598, 7105, 8288, 8359, 8623, 9139, 9799, 8568, 8760, 9626, 9078, 9050, 9048, 8988, 9138, 8871, 8971, 3930, 535, 924, 0, 824, 1965, 799, 0, 84, 0, 29, 0, 24, 0, 61, 0, 550, 1362, 454, 0, 249, 192, 0, 25, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 54, 0, 179, 0, 1620, 4085, 4298, 4573, 4116, 0, 11935, 25340, 26824, 25606, 34156, 16847, 0, 4922, 1810, 3637, 2541, 2991, 2903, 2738, 3163, 2284, 5455, 10457, 11747, 13859, 15765, 14846, 15969, 9911, 2711, 3035, 3847, 5397, 3778, 3833, 2350, 110, 73, 0, 116, 0, 945, 2919, 3127, 3363, 3312, 3636, 3551, 3065, 2977, 3229, 2442, 1143, 914, 1312, 384, 2824, 5803, 1707, 0, 101, 15, 0, 344, 0, 2817, 5650, 5195, 3303, 1321, 1171, 0, 186, 0, 45, 0, 6, 0, 0, 0, 0, 0, 0, 0, 14, 0, 96, 0, 1083, 4868, 14705, 20823, 27590, 28812, 35077, 16204, 0, 3096, 838, 2835, 1986, 2278, 1840, 1916, 1641, 2257, 1061, 3290, 0, 13299, 26777, 21372, 23219, 21704, 22303, 22015, 22105, 21998, 21839, 22757, 22551, 24667, 22359, 17801, 18606, 17119, 14991, 13905, 13506, 13973, 12440, 12020, 13701, 16724, 20942, 20481, 17873, 14164, 15778, 13158, 2572, 0, 44, 257, 1094, 958, 670, 513, 562, 533, 572, 507, 633, 249, 0, 9, 810, 1147, 170, 0, 0, 0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 33, 66, 797, 0, 4628, 15000, 18171, 20193, 21655, 22171, 23630, 26271, 27722, 28345, 26465, 22431, 18905, 15665, 7858, 2041, 2313, 1264, 120, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 28, 0, 93, 0, 817, 1960, 544, 0, 44, 0, 15, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 147, 0, 398, 0, 4756, 18869, 21236, 33035, 15747, 0, 4802, 2002, 1968, 3436, 0, 16289, 34232, 24750, 26553, 24432, 25218, 25483, 26346, 26072, 24980, 24733, 24914, 24913, 24645, 24568, 23770, 23498, 21748, 20353, 19737, 19120, 19444, 18860, 19145, 18907, 19201, 18742, 19609, 16718, 13580, 14814, 12994, 11436, 11746, 9461, 19677, 14283, 1789, 5301, 4244, 5363, 3653, 1948, 643, 0, 100, 0, 252, 775, 315, 0, 36, 0, 23, 57, 919, 1577, 2868, 2505, 1275, 1074, 132, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 36, 0, 127, 0, 1012, 2144, 1141, 361, 0, 42, 0, 12, 0, 129, 0, 623, 0, 2365, 0, 17008, 33472, 21973, 20512, 5380, 0, 4034, 5001, 7999, 8479, 13630, 10856, 3440, 2295, 0, 370, 0, 87, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 16, 0, 60, 0, 469, 1021, 862, 973, 1556, 5632, 8256, 8005, 7298, 8962, 14694, 18966, 8162, 0, 544, 0, 166, 0, 34, 0, 0, 0, 0, 0, 28856, 29099, 31053, 23348, 12547, 5093, 0, 2843, 6167, 4239, 3639, 1762, 0, 234, 0, 61, 0, 0, 26, 0, 106, 0, 1427, 6355, 8173, 7634, 8118, 7499, 8444, 6666, 13625, 28345, 28288, 35207, 15510, 0, 2790, 0, 2929, 0, 16386, 36006, 28742, 31991, 30233, 28865, 25648, 24775, 24371, 25023, 25352, 24123, 24346, 24252, 23978, 24112, 24498, 25724, 26160, 31035, 25918, 20447, 22127, 20910, 20693, 18300, 18334, 17242, 16304, 16727, 16261, 16968, 15759, 18112, 10429, 2700, 5682, 5017, 6112, 4973, 4293, 5049, 6201, 6731, 6048, 6044, 5076, 4265, 4112, 2979, 2182, 1407, 1316, 1017, 603, 297, 0, 40, 0, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 36, 0, 374, 734, 0, 1170, 4835, 5036, 10372, 15269, 17335, 23327, 25238, 36242, 16090, 0, 2740, 0, 1189, 0, 1151, 0, 2264, 0, 12845, 18464, 2359, 9860, 11109, 9167, 9987, 9153, 9133, 3748, 0, 662, 143, 273, 378, 458, 1333, 2006, 1961, 2299, 2935, 3143, 2963, 3291, 3421, 3710, 3478, 2987, 2407, 2193, 2471, 2280, 2623, 2225, 2579, 3649, 3596, 3722, 3713, 3600, 3871, 3372, 4258, 2447, 9443, 20254, 7765, 0, 1990, 0, 3548, 6589, 8265, 5330, 0, 364, 0, 102, 0, 15, 0, 0, 0, 0, 0, 0, 20, 0, 115, 0, 426, 0, 3111, 5617, 7129, 10766, 11401, 9391, 12240, 18296, 15849, 15714, 16222, 16051, 16170, 16061, 16185, 15979, 16797, 19030, 19922, 19360, 19096, 18734, 17247, 16658, 16783, 16652, 16379, 16718, 16334, 16859, 18471, 20453, 15362, 10982, 12758, 12143, 11886, 11385, 11803, 11109, 9460, 12103, 4967, 0, 135, 1212, 3994, 12488, 12128, 11484, 6734, 0, 954, 0, 265, 0, 62, 0, 45, 0, 648, 2570, 1425, 0, 348, 0, 1444, 4015, 3028, 732, 0, 63, 0, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 21, 90, 1583, 3249, 3857, 2122, 0, 8570, 16023, 14908, 16114, 16085, 16209, 15977, 16222, 14794, 16415, 6713, 0, 1282, 1361, 4525, 5240, 4625, 5096, 4191, 3809, 2714, 1467, 676, 0, 91, 0, 23, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 13, 0, 35, 0, 339, 896, 142, 99, 0, 1632, 6980, 8532, 9802, 3976, 0, 475, 0, 157, 0, 30, 0, 0, 0, 0, 0, 25, 0, 87, 0, 327, 0, 3389, 9570, 4697, 0, 17168, 26800, 21771, 26285, 26460, 27442, 27111, 28400, 29078, 29599, 30211, 29798, 30251, 30189, 30040, 29628, 29328, 26645, 24868, 24395, 22242, 20767, 19509, 18404, 18619, 18508, 17778, 17787, 17609, 17685, 17650, 17657, 17672, 17650, 17427, 15268, 13951, 14022, 13361, 15979, 18090, 18834, 19047, 21661, 22175, 24829, 15966, 2813, 2799, 2375, 1938, 1051, 1264, 1893, 1104, 0, 163, 0, 33, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 18, 0, 62, 0, 425, 490, 0, 402, 730, 639, 710, 623, 766, 334, 0, 41, 0, 7, 2, 0, 42, 0, 138, 0, 1229, 3438, 2946, 4255, 2054, 0, 219, 0, 65, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 105, 0, 392, 0, 2744, 4906, 7658, 13291, 12082, 10517, 11727, 17770, 26251, 16625, 8794, 5691, 0, 568, 0, 150, 0, 17, 0, 0, 0, 0, 0, 0, 26, 0, 137, 0, 486, 0, 3188, 3188, 0, 602, 0, 709, 0, 2031, 0, 16103, 36154, 29885, 32154, 30334, 28116, 24520, 24738, 23954, 23048, 22767, 23195, 21861, 20101, 19327, 18946, 19482, 18872, 17989, 19208, 19393, 19102, 19195, 19132, 20065, 19201, 16282, 16042, 16595, 16771, 16391, 15475, 13383, 13304, 13036, 12915, 12637, 16682, 20711, 19523, 20038, 19886, 19743, 20369, 16757, 4220, 0, 361, 0, 107, 0, 24, 0, 2, 0, 11, 0, 41, 0, 286, 403, 253, 189, 0, 29, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 12, 0, 32, 0, 290, 699, 146, 2681, 3035, 2450, 3130, 2199, 0, 7600, 18175, 18542, 23147, 22585, 22116, 22610, 22333, 20773, 23075, 21318, 22720, 26479, 25495, 25471, 26444, 24156, 29009, 12856, 0, 1606, 0, 494, 0, 370, 468, 765, 2186, 3212, 3926, 3943, 3959, 3565, 3701, 3842, 3421, 3521, 3631, 2402, 1310, 1494, 1501, 1675, 1772, 713, 0, 91, 0, 51, 0, 460, 2272, 2838, 2384, 2558, 2412, 2247, 2321, 2235, 2367, 2139, 2582, 1141, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 21, 0, 84, 0, 323, 0, 2959, 7171, 3936, 0, 9762, 23458, 26546, 31865, 31220, 32351, 31848, 31814, 31554, 31542, 30858, 31317, 27216, 23765, 24450, 23687, 24081, 23791, 24097, 23654, 24500, 21798, 19480, 19496, 19765, 18598, 19885, 7656, 0, 5888, 4600, 4801, 8831, 11410, 11593, 9863, 6943, 7427, 7076, 7340, 6835, 7387, 4570, 2370, 1530, 0, 671, 851, 668, 319, 0, 436, 170, 0, 18, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 32, 0, 106, 250, 4589, 3803, 1921, 1285, 0, 0, 4205, 18161, 24224, 26073, 25736, 26262, 24934, 24579, 22146, 17457, 18520, 16066, 18390, 12508, 764, 622, 0, 5514, 8993, 5829, 7253, 4794, 1323, 0, 122, 0, 28, 0, 6, 0, 0, 0, 0, 0, 9, 0, 44, 0, 360, 1166, 2969, 2456, 1475, 857, 0, 125, 0, 33, 0, 5, 0, 0, 0, 49, 0, 245, 0, 804, 0, 6983, 19061, 16674, 19120, 6916, 0, 2009, 0, 432, 0, 101, 0, 9, 0, 0, 0, 0, 0, 7, 0, 36, 0, 230, 0, 1785, 3256, 6455, 0, 13054, 25844, 18358, 22739, 20690, 22860, 23118, 23464, 23790, 24056, 23789, 24241, 24857, 24628, 24601, 23646, 22440, 21771, 21019, 20255, 18909, 18042, 17168, 16304, 15723, 15355, 15144, 15779, 14957, 15781, 10243, 6071, 8076, 7188, 7664, 7407, 7539, 7454, 7731, 8954, 8522, 4885, 1824, 5066, 11160, 14298, 15113, 6579, 1314, 1319, 0, 443, 423, 225, 0, 21, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 30, 0, 44, 0, 236, 1884, 0, 7959, 0, 20817, 20710, 0, 3180, 0, 890, 0, 168, 0, 1, 0, 4, 0, 4, 0, 68, 272, 0, 1417, 1150, 0, 168, 0, 48, 0, 9, 0, 0, 0, 9, 0, 48, 0, 167, 0, 1385, 3314, 2940, 3483, 3385, 3053, 3000, 2653, 2185, 2150, 723, 0, 77, 0, 70, 0, 239, 0, 815, 0, 6666, 15556, 13309, 15851, 16264, 16740, 16171, 15826, 9545, 4117, 3731, 2300, 1826, 1337, 538, 0, 59, 0, 10, 9, 0, 72, 0, 227, 0, 1888, 3129, 0, 7660, 20209, 25299, 27366, 36618, 16533, 0, 3286, 1113, 2973, 2473, 2479, 3035, 1758, 4193, 0, 15246, 31146, 25874, 28064, 26809, 27248, 26729, 26730, 26625, 26512, 26397, 26284, 25719, 26549, 26886, 21994, 19227, 19644, 19678, 19338, 18973, 19636, 19721, 19124, 19279, 19252, 19969, 20478, 20066, 22146, 23562, 27622, 15500, 1568, 2600, 1014, 1505, 2075, 1930, 2045, 1930, 2080, 1867, 2093, 177, 1444, 2778, 1340, 2304, 3605, 4156, 3449, 1646, 0, 54, 0, 16, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 55, 0, 193, 0, 1914, 6537, 8084, 8607, 8441, 9154, 8306, 13208, 17386, 14596, 15275, 6393, 0, 13998, 24967, 24366, 26922, 27649, 29564, 31047, 28810, 26203, 25073, 24454, 24935, 26503, 21046, 16939, 18014, 17694, 17465, 18377, 15940, 17578, 9804, 3457, 4436, 1047, 1909, 722, 1267, 1338, 2047, 1951, 2209, 2257, 2119, 1883, 1670, 1635, 1814, 1691, 1808, 1378, 2194, 554, 6604, 16783, 17901, 22257, 24680, 25144, 26238, 26484, 28699, 29652, 29498, 29125, 29566, 30207, 30100, 30310, 29902, 30711, 29159, 32177, 24190, 24547, 14269, 0, 1367, 0, 383, 0, 61, 0, 0, 43, 0, 184, 0, 1485, 3032, 3197, 3582, 13336, 23017, 22559, 26937, 30114, 30122, 29490, 29466, 28726, 28540, 23681, 19516, 20376, 19898, 20377, 20147, 20364, 20672, 20381, 19975, 20280, 19788, 20665, 19069, 22235, 11918, 1859, 5391, 5548, 8971, 9575, 11470, 12239, 13170, 12786, 10146, 10177, 11274, 10476, 9846, 9656, 9185, 9520, 9014, 5922, 3882, 5929, 2634, 0, 911, 406, 48, 715, 751, 231, 0, 23, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 102, 0, 766, 1520, 5454, 2491, 14238, 27776, 24455, 26614, 27091, 27383, 26684, 25824, 25126, 24963, 25564, 26227, 27665, 26415, 28588, 11283, 0, 3820, 9235, 16418, 18023, 19753, 16967, 20472, 8889, 0, 1535, 2009, 4452, 4127, 4173, 3454, 1094, 0, 126, 0, 92, 0, 217, 0, 1669, 3629, 3084, 3738, 3880, 3823, 4021, 1243, 1454, 3165, 2980, 5639, 6111, 4831, 3266, 3925, 4923, 4982, 2648, 2425, 4307, 7461, 8750, 4565, 868, 287, 527, 0, 86, 0, 21, 0, 3, 0, 0, 0, 0, 0, 7, 0, 75, 0, 323, 0, 1827, 1901, 9678, 18932, 19311, 26623, 30679, 30936, 31193, 30707, 30951, 30964, 31747, 27928, 22679, 23191, 23114, 22670, 22529, 21917, 21364, 21136, 20764, 20404, 20141, 19155, 18871, 19187, 18353, 18177, 18154, 18284, 20079, 19943, 21556, 19040, 15031, 15402, 14898, 15081, 15108, 14867, 15427, 14229, 18240, 22378, 21841, 18779, 19376, 9213, 0, 2653, 969, 1760, 621, 155, 559, 346, 341, 232, 0, 31, 0, 0, 25, 0, 197, 197, 0, 30, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 12, 0, 43, 0, 282, 282, 0, 43, 0, 12, 0, 2, 0, 0, 7, 0, 23, 0, 67, 0, 1007, 4429, 3587, 1991, 2806, 2068, 548, 0, 50, 0, 11, 0, 2, 0, 0, 0, 0, 0, 1, 0, 11, 0, 35, 27, 1410, 2809, 2644, 2069, 2157, 917, 0, 112, 0, 31, 0, 6, 0, 0, 0, 4, 0, 16, 0, 23, 153, 2625, 5617, 2096, 0, 227, 0, 69, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 182, 0, 677, 0, 12255, 22948, 27108, 28681, 35288, 17425, 0, 4997, 0, 12744, 27103, 22627, 24903, 23589, 24395, 23835, 24436, 22874, 21378, 21415, 20454, 20077, 20232, 20731, 20313, 19414, 19405, 19790, 19101, 18433, 16884, 14955, 14455, 14031, 14064, 13673, 12604, 8708, 4727, 4036, 4219, 3947, 8158, 13953, 6959, 0, 9955, 7155, 0, 1311, 588, 1455, 332, 305, 487, 0, 97, 0, 30, 19, 0, 51, 0, 680, 3212, 3410, 1295, 371, 104, 0, 13, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 72, 0, 280, 0, 1821, 2924, 4790, 4778, 0, 1286, 0, 8765, 21073, 21217, 25152, 25963, 28864, 29350, 30557, 30206, 31179, 29786, 30333, 11533, 0, 722, 958, 1674, 8826, 6107, 1014, 5480, 1520, 1094, 0, 167, 0, 27, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 50, 0, 158, 0, 1647, 6064, 7104, 9062, 7168, 12464, 19290, 19231, 21203, 22037, 24595, 27015, 19829, 4244, 0, 306, 0, 90, 0, 0, 17661, 15725, 15595, 15586, 17730, 18535, 17663, 18794, 19805, 20486, 18592, 17728, 18647, 18567, 17792, 17657, 17448, 18284, 20374, 20464, 20648, 20623, 20928, 20717, 19739, 17867, 15621, 15648, 15669, 15674, 15682, 15663, 15717, 15224, 12940, 13519, 15121, 15946, 16813, 16089, 16152, 15490, 15325, 16522, 16700, 19134, 20611, 19626, 18972, 18774, 18922, 18029, 17461, 16540, 15498, 15146, 14654, 13843, 14192, 14117, 13040, 13634, 13882, 15297, 15899, 15533, 15164, 16556, 18113, 16041, 15192, 15109, 15117, 15211, 15003, 15397, 14613, 17137, 19381, 18291, 17726, 15831, 14954, 15086, 14718, 14373, 14596, 14828, 14078, 13837, 14175, 14344, 14940, 14804, 15630, 16287, 17420, 16848, 16195, 16210, 14560, 16150, 18126, 18655, 18615, 17795, 17937, 18227, 18187, 16516, 14996, 15408, 15285, 15016, 15315, 14861, 14456, 14641, 14432, 14755, 14163, 15940, 16986, 16361, 17983, 17453, 16381, 16212, 15894, 16528, 18002, 18051, 17449, 17928, 18260, 17860, 16086, 14853, 15079, 15109, 15023, 14368, 14716, 13781, 13175, 13466, 14636, 12465, 11092, 14571, 15322, 15333, 16899, 16413, 15077, 15553, 14335, 16207, 18947, 18799, 18834, 18689, 18922, 18517, 19323, 16730, 14533, 15043, 15228, 14815, 15030, 11890, 10559, 16246, 13637, 13652, 16167, 16087, 17894, 18107, 17341, 16054, 15523, 16073, 17373, 17994, 18674, 18710, 18484, 18899, 18727, 18278, 17589, 16565, 16555, 16060, 16815, 16200, 17056, 12765, 12046, 16991, 15824, 16260, 15973, 16131, 16034, 16129, 15970, 16452, 16723, 16951, 17942, 18903, 17809, 16966, 17653, 17939, 18176, 17225, 16750, 16873, 16685, 16669, 16191, 16017, 14132, 9374, 12355, 16137, 14280, 14155, 15294, 16394, 16948, 16953, 16143, 16634, 16845, 17404, 17856, 18519, 18189, 17651, 17401, 17261, 17377, 16665, 16974, 16742, 16991, 16631, 17326, 14570, 9336, 12555, 15898, 14497, 14080, 14971, 15632, 16155, 17478, 15164, 11953, 14956, 16579, 15779, 15983, 13796, 10736, 13126, 15972, 15825, 13456, 11536, 12388, 12172, 12231, 12652, 12722, 10173, 9875, 9386, 10064, 11599, 8427, 11183, 14152, 15372, 13331, 10316, 11288, 10815, 11036, 10977, 10893, 11335, 11913, 12404, 12484, 12348, 12449, 12575, 12657, 11519, 8720, 2055, 1082, 8355, 6447, 4726, 9096, 8895, 8633, 11037, 10199, 7985, 8939, 9163, 9647, 8693, 10457, 11610, 11074, 11001, 10910, 12008, 11804, 11514, 11603, 12296, 12836, 9506, 5947, 5983, 5821, 5910, 5878, 5864, 5924, 5779, 6001, 6020, 5992, 7509, 8175, 8829, 8452, 9168, 10659, 10796, 11283, 10928, 11939, 12397, 11952, 11777, 12069, 12838, 9644, 6182, 5780, 5382, 5384, 2319, 1820, 2548, 752, 16, 1652, 4822, 5999, 6960, 7892, 8239, 8177, 7711, 8935, 10063, 9703, 9926, 9722, 9985, 9552, 10582, 9379, 7184, 6938, 5919, 5709, 4515, 2497, 3670, 6936, 3402, 0, 1501, 2429, 3586, 5786, 7034, 7201, 8599, 10439, 10003, 9996, 9766, 10753, 11286, 11272, 11409, 11166, 10695, 8912, 7445, 6441, 5437, 5829, 4367, 4057, 5811, 6221, 6549, 6408, 6518, 6392, 6586, 6208, 7570, 9784, 9877, 10010, 9699, 9792, 11003, 10503, 10128, 10393, 10472, 8649, 7156, 7757, 6568, 5310, 5593, 5596, 6014, 6273, 8196, 3129, 2554, 4459, 3052, 6706, 6218, 10505, 10880, 8777, 9620, 9421, 9864, 10362, 11345, 11300, 11440, 11677, 11709, 11771, 11617, 11928, 11343, 12484, 9174, 8546, 10998, 10044, 10874, 7446, 5689, 7850, 7467, 10065, 14572, 16852, 12513, 8795, 10025, 10053, 11314, 11591, 12106, 11813, 13643, 15431, 15391, 13924, 12211, 8348, 8127, 8018, 9163, 12159, 12795, 11803, 11515, 11275, 9048, 9771, 13936, 17640, 17137, 17488, 17255, 17457, 17205, 17643, 16265, 14905, 15636, 15514, 16222, 15949, 17124, 14451, 10791, 10941, 10599, 12315, 12633, 14168, 13385, 12557, 12205, 10777, 13817, 17191, 18361, 18865, 18049, 18742, 14542, 14229, 18462, 17154, 17176, 17267, 17091, 15930, 16024, 16042, 16875, 13530, 11048, 12389, 12121, 12287, 12248, 12173, 12384, 11916, 13719, 17329, 18508, 19510, 19656, 19987, 19303, 18080, 18421, 18418, 18232, 18186, 18227, 18773, 17776, 16062, 16460, 16794, 14313, 12356, 14343, 15251, 15340, 15747, 15653, 15504, 14212, 15295, 17007, 17691, 19562, 19340, 20904, 22954, 20329, 18690, 18708, 18618, 18691, 18661, 18658, 18695, 18607, 18812, 17894, 15042, 13062, 14456, 16066, 16012, 16749, 16421, 16860, 16136, 16238, 17659, 17773, 20827, 23144, 22561, 23895, 23027, 20199, 19188, 18953, 19309, 18860, 19056, 19331, 18001, 17192, 16642, 17074, 14944, 14805, 16469, 16248, 17568, 17757, 17421, 18429, 17866, 16409, 16800, 16778, 16465, 17234, 15606, 20707, 23848, 21601, 21822, 19262, 19022, 18879, 19090, 19092, 18012, 16349, 17649, 15466, 15154, 16834, 16003, 16765, 16825, 16084, 17610, 19624, 18988, 17424, 17327, 21090, 23044, 23781, 24919, 24982, 23651, 23527, 21296, 18999, 18888, 18722, 19055, 18747, 18465, 18007, 18151, 18104, 18077, 18194, 17951, 18316, 16831, 20243, 24083, 22272, 22385, 22432, 22957, 25080, 24570, 26456, 27519, 24526, 24260, 22080, 19918, 19044, 18853, 18999, 18784, 18917, 18238, 18259, 16968, 17881, 18299, 16819, 17720, 17520, 17239, 18739, 22190, 22942, 22385, 21132, 19438, 22761, 25709, 25599, 25832, 25557, 25961, 25279, 26606, 22297, 18056, 19149, 18653, 18614, 18355, 17451, 18019, 17965, 16704, 16709, 17328, 16808, 18324, 20751, 20335, 19350, 19157, 19807, 23148, 26326, 25912, 26002, 24951, 24142, 23643, 21125, 19125, 19385, 19127, 18966, 18980, 18668, 18902, 18009, 16791, 18071, 19095, 19244, 19246, 19205, 19289, 19133, 19484, 19177, 20852, 24784, 26543, 26638, 26768, 25832, 24231, 24166, 21982, 19684, 19608, 19510, 19430, 19507, 19149, 19096, 18880, 16122, 17513, 18506, 17989, 18636, 17527, 19078, 22144, 21997, 19725, 20025, 19100, 22899, 26968, 26849, 27037, 25104, 24441, 25004, 22431, 20616, 21097, 20899, 20927, 21093, 20269, 19066, 19056, 20063, 18807, 22369, 25496, 22739, 22695, 25297, 26140, 26427, 22629, 19668, 24863, 26755, 26952, 26961, 26612, 25359, 24949, 22783, 20002, 19885, 19403, 19671, 19770, 19112, 18921, 19170, 19706, 19179, 21323, 25884, 26103, 25294, 26116, 26817, 27290, 27411, 27499, 27251, 27749, 26772, 29408, 28304, 25146, 26328, 24538, 25147, 21881, 19510, 20200, 21501, 24315, 21865, 19969, 19362, 20950, 25639, 27324, 27437, 27484, 27601, 27965, 28238, 28478, 28081, 28151, 28098, 28233, 26880, 29660, 29712, 26039, 25451, 25264, 22238, 19112, 19999, 19502, 19309, 18987, 19049, 18968, 19090, 18883, 19287, 18005, 17039, 18474, 18851, 22112, 22478, 20050, 17525, 17722, 24204, 27017, 26791, 25880, 24219, 24608, 21842, 19806, 18700, 17861, 19261, 19147, 19420, 19095, 18009, 15588, 17513, 19489, 18653, 17683, 17478, 18075, 18603, 20385, 19722, 16953, 15457, 17433, 19931, 20526, 20435, 20442, 20490, 20368, 20641, 19678, 18420, 18752, 18834, 17677, 17198, 19020, 16953, 17092, 19701, 19604, 18769, 17642, 19082, 20377, 21924, 22742, 21698, 19500, 23327, 27540, 25667, 25105, 24556, 24317, 23902, 24084, 24188, 23032, 23023, 23689, 24100, 23835, 23043, 19444, 18863, 18075, 21784, 26130, 24745, 25463, 25042, 25324, 25061, 25772, 26804, 25668, 27709, 29362, 29309, 26661, 23666, 23806, 23754, 23854, 22564, 22511, 23923, 23204, 23110, 19898, 17227, 18327, 17997, 18329, 21478, 24697, 23595, 23680, 24984, 25244, 24953, 23994, 23626, 23750, 25370, 28677, 25669, 21527, 21587, 21798, 22337, 22436, 22475, 22360, 22596, 22142, 23067, 20051, 17177, 17720, 17485, 17938, 18573, 18294, 18552, 22271, 22864, 22467, 21320, 19903, 21665, 21879, 21863, 19429, 16720, 17274, 17528, 18698, 19278, 18521, 18617, 19189, 18719, 17531, 17245, 17315, 16741, 16582, 17021, 17119, 17908, 17211, 19252, 22273, 21570, 21602, 21589, 21464, 21783, 21162, 22359, 19125, 21158, 27814, 24011, 20268, 20786, 22521, 21801, 21373, 18351, 15789, 15883, 15722, 15133, 14863, 15851, 18196, 19078, 20218, 21784, 20405, 20759, 19187, 24178, 29283, 27836, 27762, 22218, 22604, 25921, 26182, 25239, 23265, 26064, 29893, 25162, 19367, 17073, 15063, 15691, 15439, 15464, 15647, 15093, 17844, 26145, 29339, 28437, 28856, 28202, 28359, 28961, 28691, 26933, 23447, 23657, 25540, 25421, 25434, 26375, 26518, 26782, 29310, 23475, 17268, 18227, 17914, 19229, 19475, 18896, 24243, 27758, 27348, 28868, 29257, 29043, 29140, 29526, 29765, 29993, 30238, 29693, 29363, 29449, 29403, 29449, 29375, 29496, 29475, 30409, 24958, 20731, 21423, 20040, 20325, 20326, 24815, 27556, 26779, 28459, 29334, 30063, 30799, 30426, 30295, 30600, 30871, 31072, 31054, 30491, 29852, 29885, 29944, 29881, 30215, 30821, 30979, 31118, 29744, 27974, 27288, 27140, 27266, 27775, 29311, 30105, 30071, 30097, 30106, 30057, 30166, 29936, 30728, 31734, 31748, 31865, 31616, 31344, 31351, 31288, 30969, 31511, 31600, 31587, 31369, 26871, 24729, 24047, 23613, 23778, 26473, 29175, 29300, 30061, 29687, 30650, 30795, 30179, 29301, 30055, 30792, 31121, 31603, 31488, 31372, 31251, 31422, 31359, 31613, 32157, 32283, 32291, 32238, 32348, 32141, 32566, 31056, 29120, 30341, 30658, 30015, 30720, 30616, 29886, 30137, 29832, 29138, 30318, 31421, 31230, 31579, 31798, 31496, 31241, 31855, 32337, 30837, 30789, 31125, 31246, 28064, 25069, 26031, 24977, 27179, 29702, 30492, 30227, 29457, 30092, 30220, 30301, 30890, 30605, 29946, 30436, 29719, 30886, 28882, 32924, 17311, 0, 18601, 34811, 29227, 32526, 30837, 30147, 27861, 27572, 27442, 28841, 31138, 31696, 31644, 30977, 30716, 30394, 30729, 30795, 29844, 30035, 28940, 33094, 29409, 38629, 12229, 12006, 38471, 29030, 31412, 26864, 27758, 27115, 28039, 27805, 27583, 27396, 27220, 27272, 27261, 27237, 27306, 27151, 27600, 27713, 27961, 27444, 26860, 26986, 28462, 31555, 31908, 32914, 30885, 28635, 29052, 28688, 27924, 26676, 26936, 27329, 27261, 26958, 26663, 26477, 26782, 26952, 30449, 30469, 28185, 28001, 27063, 27881, 28099, 27850, 27295, 27355, 27464, 27916, 30397, 30475, 29516, 29888, 29607, 29922, 29458, 30305, 27638, 25339, 26565, 25519, 25439, 25394, 26080, 27212, 27733, 27818, 27594, 27082, 26945, 27749, 27531, 26825, 26682, 26630, 27372, 28226, 28504, 28328, 28042, 27847, 27253, 27162, 23580, 19616, 20991, 22787, 22944, 23286, 23919, 24133, 24655, 25359, 26761, 27293, 26974, 27112, 27022, 27105, 26996, 27182, 26709, 27025, 27872, 28549, 28277, 27102, 27373, 26447, 26153, 22725, 18193, 19145, 20575, 20850, 22175, 21845, 21594, 22385, 24781, 25826, 25130, 26010, 25111, 24428, 25235, 25819, 25831, 25574, 25045, 25640, 26273, 26587, 26825, 25834, 25268, 24503, 24014, 21904, 20115, 20686, 20340, 20638, 20281, 20842, 19508, 21200, 25017, 22446, 23049, 24187, 23114, 23996, 24070, 24468, 23430, 24113, 25210, 24733, 25633, 25597, 25599, 24314, 24581, 23146, 18976, 17817, 17174, 18100, 19332, 18639, 18153, 16947, 16654, 20672, 24490, 23451, 22665, 22906, 21478, 22799, 23760, 23164, 23313, 23230, 23239, 23318, 23114, 23535, 22505, 23084, 20666, 17706, 16878, 16717, 17395, 16961, 16524, 17033, 14553, 14788, 18635, 19867, 20069, 19461, 20564, 19772, 21986, 22740, 21920, 21055, 22220, 23386, 22582, 24527, 23539, 22736, 22169, 21820, 19983, 17795, 16800, 16335, 17672, 17845, 17111, 16786, 17219, 17138, 17039, 17351, 16649, 19042, 22073, 23376, 23106, 21235, 22138, 22305, 21643, 22639, 24158, 22785, 21817, 20856, 20865, 19634, 17886, 17171, 16486, 17686, 17780, 17762, 19676, 15520, 15266, 19532, 20745, 20206, 20560, 21945, 21759, 23847, 23164, 21242, 21470, 22518, 21871, 23148, 23408, 22073, 22083, 21906, 22176, 21726, 22587, 19844, 17333, 18362, 18581, 19816, 16193, 16594, 19428, 20379, 20656, 21056, 22518, 22139, 22839, 22693, 22012, 21329, 21725, 21178, 22637, 23224, 21837, 21203, 20434, 19510, 18148, 17986, 17428, 17429, 17617, 18037, 17684, 18792, 15794, 15922, 19556, 19534, 19990, 21269, 22661, 22196, 22483, 22222, 22582, 21682, 21727, 22979, 23553, 23490, 21800, 21984, 20861, 18916, 17957, 17781, 17661, 16836, 17666, 18361, 18752, 18170, 18248, 19715, 19598, 19006, 20929, 21741, 21440, 22309, 21499, 21584, 21494, 21772, 21674, 22695, 23571, 21933, 21404, 20919, 19499, 17967, 17458, 17215, 17276, 17274, 17219, 17356, 17063, 17941, 18362, 19141, 19468, 20840, 20952, 21250, 21650, 20223, 20671, 20096, 21659, 21759, 21424, 22393, 21239, 20858, 19144, 18110, 18092, 17025, 17117, 17507, 17342, 18234, 16630, 13878, 14024, 16866, 20497, 19032, 18687, 20869, 21528, 21711, 21016, 20319, 21407, 21918, 21841, 21801, 21957, 21622, 22317, 20049, 17987, 18406, 17358, 17611, 17983, 17725, 18516, 18456, 14876, 15903, 19418, 19824, 17425, 18205, 21005, 21556, 21166, 20552, 20271, 21226, 22648, 22066, 21680, 22257, 22211, 20969, 20656, 18920, 17502, 17623, 17279, 17508, 17597, 17339, 18487, 16501, 14669, 15270, 14932, 15193, 14916, 15307, 14582, 17136, 20813, 19559, 20336, 21661, 21259, 21296, 22314, 20481, 18618, 18434, 17369, 18019, 17068, 16943, 18018, 16850, 17664, 14332, 12541, 14264, 15704, 19316, 17319, 15437, 18056, 19659, 19649, 18956, 18692, 20847, 21181, 21270, 21778, 21343, 21993, 21505, 20166, 19731, 19854, 19742, 19889, 19660, 20128, 17942, 11972, 12807, 14282, 15933, 19078, 17108, 16671, 18298, 19762, 19283, 18344, 20324, 21370, 21545, 21732, 21596, 22202, 22078, 21408, 21297, 19279, 17791, 18005, 17573, 17992, 18133, 18303, 18343, 15975, 14197, 16855, 19065, 19490, 17907, 18692, 21902, 22765, 23037, 22947, 22996, 22957, 23005, 22935, 22971, 21980, 21994, 22588, 19873, 18501, 18416, 17879, 18036, 18401, 18253, 19890, 16855, 16778, 19727, 19901, 19961, 18335, 20744, 23043, 22191, 22506, 22895, 22784, 24197, 23433, 24043, 24299, 23155, 22877, 22761, 22957, 22107, 19770, 18343, 18544, 18502, 19740, 20637, 20375, 20510, 20434, 20477, 20441, 20720, 22521, 24045, 25279, 24644, 23290, 24358, 24805, 24150, 24208, 24219, 23799, 23222, 23110, 23334, 22336, 19867, 18210, 18467, 18482, 19270, 20083, 19928, 19962, 20907, 22374, 23601, 23725, 23859, 24519, 24845, 25263, 25425, 25145, 25257, 25030, 25101, 25379, 25165, 25291, 25160, 25351, 25029, 25647, 23688, 22059, 23166, 23138, 23446, 20872, 20588, 22987, 24002, 24218, 24986, 25048, 24599, 25665, 25800, 25665, 25891, 25720, 25026, 25733, 26364, 25557, 25105, 23659, 23332, 23155, 23165, 22407, 21338, 21993, 22488, 23177, 23715, 22372, 22451, 24705, 23855, 24744, 25893, 25524, 25735, 25583, 25726, 25523, 26196, 27202, 26229, 25630, 25467, 25080, 24199, 24495, 24466, 22987, 20521, 19714, 19135, 20489, 22266, 20881, 19939, 19562, 22446, 23524, 23976, 25138, 25618, 25701, 26339, 26330, 26510, 26728, 26053, 25797, 25065, 26025, 25062, 24314, 24052, 23644, 23768, 23768, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 886, 0, 3148, 0, 20631, 20631, 0, 3148, 0, 886, 0, 170, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 28, 28, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 3, 0, 34, 167, 310, 463, 187, 0, 20, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 18, 0, 120, 113, 0, 24, 0, 0, 82, 272, 410, 310, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 10, 230, 234, 285, 193, 0, 20, 66, 402, 405, 348, 409, 505, 322, 69, 54, 0, 14, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 16, 68, 10, 123, 87, 0, 0, 129, 458, 406, 555, 714, 515, 440, 459, 441, 468, 422, 510, 225, 0, 28, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 7, 0, 69, 190, 44, 108, 94, 0, 14, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 40, 83, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 24, 0, 161, 161, 0, 24, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 78, 78, 0, 12, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 0, 100, 100, 0, 15, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 882, 0, 3131, 0, 20565, 20876, 0, 3204, 0, 885, 0, 171, 0, 0, 0, 0, 0, 0, 3, 0, 12, 0, 236, 170, 0, 24, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 39, 39, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 39, 0, 277, 481, 608, 688, 419, 774, 892, 289, 0, 28, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 97, 0, 344, 0, 2299, 2587, 0, 895, 225, 654, 770, 360, 92, 25, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 171, 0, 958, 0, 3265, 0, 20875, 20678, 0, 3133, 0, 853, 0, 304, 0, 20, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 10, 0, 70, 58, 0, 0, 99, 192, 155, 367, 365, 142, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 9, 0, 104, 300, 113, 307, 221, 0, 32, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 21, 0, 141, 141, 0, 21, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 9, 0, 64, 64, 0, 9, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 17, 17, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0);

--  Datos de 17 a 32
--    type t_reg_datos is array (0 to 32783) of integer range 0 to 30000;
--    signal reg_datos_debug : t_reg_datos := (0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7398, 0, 926, 0, 275, 36, 2031, 2839, 1243, 553, 213, 0, 29, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 37, 0, 131, 0, 1059, 2378, 2000, 2145, 2145, 2000, 2378, 1059, 0, 131, 0, 37, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 343, 3172, 6075, 6687, 7011, 7447, 7786, 8077, 7321, 6657, 6927, 6651, 7053, 6372, 7693, 3400, 0, 422, 0, 120, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 18, 0, 53, 72, 2330, 4330, 4188, 4703, 5096, 5148, 4899, 5932, 6276, 5573, 5720, 5719, 5694, 6447, 6891, 6848, 6726, 7045, 6408, 7710, 3414, 0, 418, 0, 100, 0, 0, 106, 0, 1281, 4661, 5239, 4820, 4923, 4231, 4029, 4218, 4406, 4064, 2687, 759, 0, 76, 0, 20, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 43, 0, 150, 0, 1271, 3189, 3013, 3845, 4313, 4584, 4374, 4104, 3925, 4034, 3337, 5464, 8372, 8383, 8792, 9127, 7974, 7619, 7771, 7794, 7669, 7944, 8916, 10542, 7549, 4090, 4229, 3070, 2688, 1854, 1569, 1427, 1031, 257, 0, 22, 0, 2, 0, 0, 21, 0, 77, 0, 856, 3293, 4093, 4150, 4234, 3724, 1142, 0, 117, 0, 33, 0, 17, 0, 50, 0, 180, 0, 1713, 5376, 6789, 7431, 8472, 8908, 9190, 10573, 10186, 9869, 8011, 7106, 5630, 4477, 7359, 9334, 9561, 9228, 7426, 6264, 6607, 6393, 6599, 6323, 6770, 5916, 8670, 11311, 10374, 10968, 9376, 8148, 7941, 7863, 8025, 8014, 6970, 6742, 2547, 0, 296, 0, 84, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 165, 0, 576, 0, 4707, 10834, 8387, 8532, 8500, 9135, 9318, 9168, 8999, 9673, 9480, 9222, 9262, 8493, 7765, 6444, 4886, 4183, 1877, 1676, 4262, 4737, 6244, 7660, 7449, 7589, 7787, 7718, 7276, 7167, 7155, 7278, 6979, 6755, 7079, 6763, 7239, 5306, 3566, 4121, 3787, 4059, 3755, 4268, 2296, 0, 3125, 7445, 7848, 8490, 8494, 5397, 803, 0, 28, 0, 8, 0, 0, 0, 0, 22, 0, 74, 0, 1293, 6945, 10058, 10187, 10141, 11116, 11857, 11743, 12397, 13062, 13261, 12281, 10072, 9394, 10037, 8406, 7201, 7212, 7004, 7390, 6693, 8072, 3569, 0, 443, 0, 126, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 41, 0, 244, 753, 4318, 7913, 7977, 7688, 7043, 7270, 5479, 2137, 389, 0, 31, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 201, 1161, 2548, 3124, 3213, 2955, 3871, 6994, 7591, 5986, 5644, 5470, 5176, 5166, 5285, 5345, 5059, 5282, 4961, 4750, 4911, 4652, 2360, 50, 59, 0, 18, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 19, 0, 65, 0, 507, 943, 147, 0, 0, 0, 0, 13, 0, 80, 0, 284, 0, 3234, 7798, 8202, 8966, 9303, 9929, 10544, 11395, 11752, 12013, 11894, 12019, 11829, 12159, 11519, 13446, 14416, 13801, 14842, 15125, 15452, 15597, 15577, 14611, 13806, 13101, 12713, 12136, 11530, 10066, 8829, 6768, 2378, 1903, 3409, 4879, 6814, 9855, 12785, 14234, 15494, 16190, 17317, 17561, 17771, 17966, 16769, 13675, 7306, 2259, 558, 0, 54, 0, 0, 91, 0, 356, 0, 2888, 6531, 4711, 4553, 3570, 4190, 3425, 2164, 4656, 4482, 3055, 3382, 6442, 8043, 6555, 5471, 4700, 5212, 5409, 6221, 7016, 7497, 8041, 8666, 9385, 9755, 10329, 10958, 11043, 11579, 11797, 11808, 11343, 10734, 10066, 10164, 14329, 15505, 14276, 14746, 14483, 14655, 14514, 14686, 14262, 14188, 14640, 14177, 13960, 13648, 13662, 13128, 12597, 11381, 10920, 4054, 0, 443, 0, 45, 289, 1072, 1369, 2283, 3266, 3837, 3517, 1099, 0, 220, 0, 420, 0, 3285, 8322, 8135, 8984, 9151, 9923, 9486, 9673, 10470, 10485, 10596, 10397, 10751, 10109, 11405, 6843, 217, 161, 0, 30, 8, 0, 1093, 3193, 4462, 5211, 5487, 5807, 6242, 6318, 6800, 7446, 7764, 7818, 8431, 9324, 10029, 10071, 9460, 9558, 9565, 9275, 9040, 9053, 9240, 9399, 9180, 8075, 6972, 3304, 118, 63, 0, 21, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 7, 122, 160, 0, 159, 0, 506, 0, 3273, 7938, 7827, 8926, 8919, 9333, 9263, 9377, 9346, 9312, 9432, 9538, 9564, 9015, 7979, 7478, 7669, 7458, 7789, 7213, 8319, 5023, 3741, 6476, 6714, 8869, 7261, 6612, 7187, 9271, 8286, 7330, 9470, 9842, 10604, 10494, 10030, 9890, 9322, 6839, 1935, 0, 191, 0, 53, 0, 1, 9, 0, 84, 0, 296, 0, 2727, 7743, 8841, 10081, 10379, 10831, 10869, 10895, 10835, 10955, 10711, 11220, 9455, 6382, 3403, 4465, 7781, 8695, 9631, 9715, 10080, 10550, 10754, 10682, 10836, 10815, 10464, 10559, 9560, 8467, 3020, 0, 342, 0, 97, 0, 15, 0, 0, 15, 0, 54, 0, 817, 4020, 6100, 6732, 7521, 7899, 8425, 8750, 8673, 8680, 8731, 8599, 8883, 7941, 6998, 6899, 5984, 5586, 5777, 5689, 5858, 6399, 6485, 6532, 6499, 6734, 6584, 6740, 5546, 4569, 5102, 5436, 6424, 7413, 7261, 7103, 7319, 7032, 7656, 7358, 7480, 8188, 7169, 7297, 7096, 6758, 6594, 5202, 1597, 0, 164, 0, 46, 0, 5, 0, 0, 37, 0, 138, 0, 1141, 3095, 4948, 6878, 6935, 6212, 5460, 1927, 0, 152, 11, 0, 667, 194, 2926, 7105, 8876, 4773, 0, 674, 0, 2993, 7109, 6541, 7088, 6650, 6535, 6339, 6658, 6021, 6984, 3002, 0, 353, 0, 21, 104, 0, 547, 0, 4624, 11208, 9548, 9367, 8274, 8598, 8067, 11709, 14305, 14374, 12749, 12611, 11179, 6784, 6476, 6412, 6346, 6110, 5701, 5505, 4447, 4653, 5933, 7512, 9394, 10053, 11358, 13371, 14801, 14927, 15033, 14886, 15178, 15094, 15129, 14588, 13639, 13635, 13641, 13798, 13438, 14140, 12829, 15455, 6839, 0, 849, 0, 243, 0, 50, 0, 6, 0, 22, 0, 166, 304, 178, 74, 0, 0, 73, 82, 0, 12, 0, 3, 0, 1, 0, 7, 0, 32, 0, 440, 2287, 4673, 6314, 6653, 6719, 6877, 6931, 6922, 6920, 6930, 6904, 6959, 6773, 6453, 5829, 5485, 5611, 6053, 6592, 6865, 7081, 7191, 7583, 7876, 8189, 8514, 8990, 9409, 9391, 9653, 9895, 10050, 10277, 8951, 9562, 4793, 908, 1754, 4199, 7542, 7568, 8262, 7842, 7690, 3879, 3623, 6981, 7658, 8194, 8616, 8979, 8955, 8797, 9187, 8420, 9950, 5327, 3658, 8167, 9641, 11989, 12236, 12846, 12874, 12758, 12983, 8859, 5953, 6871, 6464, 6816, 6588, 6645, 6645, 6803, 6802, 6624, 5967, 3647, 1341, 3619, 6508, 6397, 6680, 6935, 7054, 7362, 7400, 7572, 7382, 7203, 7495, 7294, 7275, 7401, 7339, 7396, 7333, 7414, 7257, 8044, 9806, 2975, 105, 0, 2997, 0, 20866, 20097, 0, 5661, 5563, 14788, 13963, 15950, 15943, 16175, 16345, 16331, 16376, 16133, 16259, 13668, 11685, 12316, 12176, 12555, 12427, 12567, 12525, 12872, 13106, 13248, 13480, 13537, 13838, 13948, 13762, 13721, 13747, 13680, 13819, 13615, 13069, 4422, 0, 478, 0, 140, 0, 65, 121, 116, 211, 600, 3904, 7859, 6747, 10520, 13979, 14173, 12311, 9600, 10658, 9060, 9454, 3522, 0, 20, 963, 2050, 8002, 14387, 13876, 15165, 13975, 9688, 7512, 8564, 8594, 8621, 8466, 8398, 8420, 8402, 8425, 8393, 8462, 8392, 8462, 8705, 9105, 9337, 9191, 9322, 9543, 9534, 9632, 8955, 7489, 5424, 4365, 4210, 4296, 4876, 4851, 6195, 7253, 8048, 8197, 7464, 6641, 1989, 0, 200, 0, 52, 0, 0, 58, 0, 230, 0, 1926, 4809, 4816, 5331, 5153, 5176, 5291, 4968, 6167, 7883, 8041, 8070, 8133, 8494, 8777, 8295, 8762, 7020, 9903, 13372, 12161, 12925, 11032, 10216, 10380, 10511, 10369, 11418, 13554, 14177, 14493, 14597, 14365, 13783, 13496, 13443, 13308, 12975, 13013, 12882, 12983, 11857, 9742, 9315, 9572, 9870, 9978, 9902, 10012, 9853, 10099, 9590, 12161, 17848, 6718, 0, 734, 0, 143, 500, 3754, 5329, 5690, 6270, 6425, 6856, 6813, 7009, 6911, 6911, 6483, 5445, 2630, 0, 4494, 10005, 9117, 10045, 9832, 10090, 9955, 9820, 9993, 9833, 9868, 9992, 9963, 10248, 10204, 9957, 9858, 9888, 9870, 9879, 9887, 9861, 9732, 8767, 10492, 7682, 4340, 4484, 4158, 4214, 3808, 4772, 5298, 6393, 6537, 6413, 6674, 6679, 6317, 6250, 6264, 5143, 5166, 5473, 5564, 4628, 3848, 4015, 4952, 6299, 6159, 6626, 5702, 5561, 2616, 390, 955, 624, 853, 576, 791, 704, 741, 733, 722, 756, 618, 353, 301, 33, 62, 0, 861, 3253, 4386, 4275, 4992, 2013, 0, 202, 0, 0, 2196, 9547, 12916, 13723, 15022, 14890, 16758, 17778, 17724, 17915, 18289, 18102, 16803, 16141, 14786, 14205, 13107, 14858, 7646, 860, 2865, 1765, 2272, 2025, 2087, 2171, 1932, 2432, 900, 518, 3496, 4036, 4237, 6112, 7343, 7623, 8135, 8233, 8392, 8583, 8693, 8514, 7659, 8242, 3184, 0, 389, 0, 547, 2329, 2792, 231, 1015, 2698, 2539, 2410, 1225, 284, 0, 97, 0, 277, 0, 2300, 6080, 7331, 8531, 8191, 8228, 8454, 7885, 9087, 5308, 3138, 5837, 5351, 5874, 6145, 6528, 6720, 7204, 7034, 7508, 6609, 6652, 2740, 0, 333, 0, 94, 0, 18, 0, 0, 0, 0, 0, 10, 0, 51, 0, 174, 0, 1633, 4944, 5391, 6519, 6985, 7257, 8070, 8199, 8220, 8153, 8293, 8013, 8564, 7174, 7308, 3253, 0, 410, 0, 115, 0, 29, 0, 31, 0, 130, 0, 1332, 5179, 6519, 6817, 7711, 8033, 7953, 8323, 8448, 8608, 8746, 8687, 8787, 8865, 7870, 6298, 1770, 136, 1629, 1151, 1439, 1329, 1279, 1232, 1268, 1272, 1243, 1306, 1186, 1428, 632, 0, 78, 0, 22, 0, 4, 0, 18, 0, 90, 0, 320, 0, 2743, 7343, 8195, 9804, 10185, 11092, 11752, 10766, 14488, 17847, 17665, 17899, 18381, 14998, 11867, 12476, 11875, 12221, 11884, 11818, 11954, 11872, 11802, 12032, 12049, 12083, 12006, 12161, 11868, 12417, 11245, 14430, 18691, 18330, 18733, 18082, 17412, 14439, 12597, 13482, 13172, 13116, 13092, 12357, 12266, 11789, 11489, 11452, 11411, 11302, 10995, 8980, 7650, 2835, 0, 330, 0, 93, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 162, 0, 569, 0, 4560, 10247, 8738, 9800, 9259, 9594, 9592, 9534, 9551, 9638, 9434, 9322, 8825, 7551, 6451, 6029, 5961, 5273, 5115, 5731, 6250, 6522, 7201, 8167, 9003, 9758, 9704, 9900, 9943, 10089, 9572, 8970, 9095, 8921, 8888, 9232, 9252, 9087, 9087, 9179, 8947, 9411, 8539, 10287, 4551, 0, 565, 0, 161, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 514, 4272, 8918, 9806, 9963, 10639, 11334, 11244, 11529, 11786, 11924, 11147, 14301, 18201, 18119, 18601, 18768, 19003, 18681, 18878, 18640, 19025, 18337, 19698, 15267, 10870, 11824, 11369, 9952, 7747, 7719, 7541, 7771, 7554, 6760, 7245, 4535, 0, 5335, 12919, 12805, 14590, 12112, 10436, 3865, 0, 523, 0, 356, 0, 1992, 5398, 5486, 6534, 6466, 7150, 2824, 0, 335, 0, 96, 0, 35, 0, 79, 0, 277, 0, 2481, 7088, 7760, 8263, 8340, 8777, 8686, 8712, 8871, 8911, 9052, 8809, 8546, 8837, 9277, 9158, 9547, 10269, 10297, 10079, 9104, 8827, 8838, 8571, 8120, 7189, 5538, 1514, 0, 143, 0, 50, 0, 52, 0, 153, 0, 1240, 2792, 2335, 2533, 2481, 2406, 2661, 1696, 411, 282, 582, 1012, 993, 970, 1094, 1138, 937, 806, 865, 793, 1434, 622, 3565, 6967, 6752, 7851, 7231, 7277, 7005, 7250, 7236, 8510, 3526, 0, 481, 63, 1320, 819, 840, 690, 179, 216, 311, 221, 10, 33, 0, 174, 0, 577, 0, 4801, 11806, 9114, 11596, 4707, 0, 567, 0, 172, 0, 34, 0, 0, 0, 12, 0, 58, 0, 204, 0, 1833, 5019, 5266, 6208, 6608, 7142, 7665, 7980, 8234, 8106, 8357, 8466, 8959, 10017, 10701, 11472, 11797, 11836, 11896, 11849, 11914, 11805, 12013, 11348, 10871, 11748, 12406, 12488, 12093, 12456, 12860, 13067, 14144, 14641, 14245, 14223, 14238, 12501, 11399, 6689, 702, 0, 0, 7, 0, 0, 0, 67, 58, 179, 143, 113, 294, 442, 607, 671, 747, 1003, 397, 0, 128, 0, 26, 0, 6, 0, 0, 0, 0, 14, 0, 75, 0, 268, 0, 2429, 5173, 4801, 4349, 3616, 1583, 0, 198, 0, 53, 0, 10, 0, 0, 0, 4, 0, 17, 0, 56, 0, 678, 2704, 3207, 3806, 4825, 5698, 6416, 6666, 6386, 4544, 3651, 3955, 3678, 4056, 3379, 5544, 7924, 7527, 8162, 8327, 8874, 9498, 10123, 10521, 11130, 11086, 11757, 10416, 10463, 5469, 760, 2304, 1524, 1834, 1803, 1778, 1596, 1560, 1454, 1390, 1401, 1500, 1538, 1634, 1604, 1584, 1520, 1488, 1496, 1518, 1556, 1508, 1526, 1534, 1549, 1510, 1588, 1441, 1736, 765, 0, 73, 0, 0, 151, 0, 1156, 1115, 0, 232, 0, 56, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 64, 64, 29288, 29190, 29799, 29660, 29971, 29658, 29593, 29474, 29740, 29229, 30313, 26018, 16918, 13316, 10022, 4015, 2367, 718, 7313, 16896, 19284, 25190, 27309, 28028, 29280, 29731, 30547, 30663, 30485, 30130, 29103, 27038, 26930, 28102, 28147, 28371, 26908, 28585, 24841, 19186, 14137, 8677, 5425, 1323, 2633, 715, 6246, 13540, 13922, 19587, 22084, 21630, 21618, 22031, 20957, 24697, 28095, 26724, 28751, 28554, 29091, 30145, 30081, 30273, 28282, 28463, 27689, 20897, 14809, 10398, 4889, 2961, 4284, 2343, 6299, 12893, 14951, 21122, 24639, 25467, 27315, 28169, 29180, 29261, 30119, 30674, 30957, 31307, 31015, 31155, 31138, 31477, 30471, 29014, 29591, 28742, 30177, 27594, 32694, 16409, 1706, 4526, 6536, 15707, 18069, 22474, 23414, 25137, 27401, 28510, 29642, 30890, 30211, 30526, 30526, 30087, 30450, 30164, 30180, 29995, 29180, 28383, 30227, 26113, 20894, 20563, 12961, 5360, 3789, 4287, 2621, 7609, 14835, 21007, 26847, 28180, 27999, 26803, 27174, 27068, 26983, 27274, 26606, 28909, 31601, 31352, 30346, 28858, 29040, 30583, 26564, 21769, 18386, 11597, 5847, 4357, 4468, 4261, 2667, 7640, 16310, 20094, 23771, 25890, 27809, 29780, 30946, 31495, 31764, 31510, 31001, 30610, 31583, 31501, 31060, 30516, 29956, 31166, 28112, 21443, 16549, 14895, 15310, 15110, 15217, 15163, 15189, 15096, 15781, 22143, 27991, 29187, 30391, 31648, 32714, 32532, 32608, 32401, 31233, 31374, 31813, 30924, 30566, 28458, 28762, 26247, 18588, 15293, 11585, 8309, 5609, 5634, 5173, 4234, 2180, 8558, 15317, 16501, 23255, 23391, 26471, 30288, 31284, 32227, 31669, 32013, 31847, 31941, 31877, 31930, 31890, 31680, 27829, 18659, 15382, 12163, 7922, 5807, 5419, 4571, 4117, 1633, 7707, 14471, 15136, 22646, 23773, 24980, 28663, 30392, 29903, 29978, 30003, 29419, 29007, 29065, 28177, 26992, 24517, 22007, 22571, 17351, 11512, 10643, 6667, 3878, 4338, 3968, 3157, 3016, 2779, 3376, 2207, 4386, 14, 14632, 30945, 27073, 29243, 28596, 29340, 29346, 28769, 27269, 23973, 21034, 19834, 17787, 14302, 10282, 8647, 5774, 3717, 4577, 4289, 3253, 3080, 260, 6790, 13921, 13034, 15603, 15751, 20972, 27698, 27525, 28134, 29825, 29136, 28839, 26932, 24179, 17606, 14008, 15103, 14359, 15136, 14031, 16034, 9632, 3242, 4988, 3296, 2257, 2203, 1394, 7765, 13260, 13601, 13130, 18318, 30516, 26940, 25458, 29623, 29484, 31219, 25887, 17213, 14363, 14494, 14842, 12454, 9054, 5460, 3460, 4163, 3762, 3295, 3633, 3011, 2905, 833, 5556, 12052, 12102, 13162, 13366, 13141, 13673, 12630, 14561, 10774, 22509, 28519, 15034, 14846, 14360, 13490, 8242, 3124, 3003, 3263, 3507, 3456, 2955, 2838, 2359, 3441, 1041, 6633, 12660, 9689, 13484, 10446, 22255, 31608, 28779, 32108, 30385, 30569, 32195, 25007, 17612, 20130, 17531, 11746, 6880, 3095, 2475, 2992, 2843, 2846, 2997, 2597, 3429, 1706, 7027, 10692, 11899, 10343, 21138, 32719, 29215, 31825, 30174, 31526, 31840, 30921, 25038, 20453, 20429, 15106, 10442, 6582, 2675, 2149, 3181, 3140, 2641, 2699, 2958, 3544, 1732, 6877, 10721, 11350, 9952, 21371, 34273, 30378, 33474, 29669, 36473, 16577, 0, 2420, 0, 799, 568, 0, 3312, 4446, 1926, 3325, 2764, 3094, 2772, 4480, 2464, 6664, 13722, 10569, 15675, 19299, 29028, 29045, 38219, 11198, 15235, 24986, 0, 20141, 33050, 26577, 28830, 25237, 23333, 17336, 10296, 4437, 2194, 3509, 3000, 3462, 3478, 4554, 2501, 8253, 13613, 12119, 12598, 12866, 11684, 14442, 6117, 1536, 0, 16380, 37339, 29279, 31242, 29955, 29303, 24793, 21231, 13305, 4058, 2772, 3015, 3411, 3064, 4864, 2475, 7650, 14033, 17494, 27307, 21216, 32159, 17034, 0, 3827, 0, 3579, 0, 16516, 37098, 29538, 31779, 29978, 29912, 25741, 22828, 23911, 22946, 24181, 22206, 25966, 13707, 1070, 9993, 15088, 25013, 22463, 30335, 14754, 0, 955, 3273, 0, 22812, 16523, 10027, 40248, 27990, 32819, 28927, 29529, 25939, 18545, 8945, 2640, 3059, 4031, 3272, 4386, 2235, 7529, 13397, 16940, 26179, 27372, 23918, 35354, 16587, 0, 2543, 0, 1565, 0, 2526, 0, 16175, 34684, 27516, 25923, 20509, 13748, 3137, 2969, 3870, 3376, 3820, 4000, 9662, 13334, 20153, 30355, 21616, 31557, 16655, 0, 3418, 0, 3445, 0, 16429, 36916, 30452, 32567, 30394, 31279, 28478, 25517, 15658, 6865, 4261, 2908, 4684, 4078, 3592, 3263, 4338, 2066, 6425, 0, 22004, 20096, 0, 3641, 0, 1337, 803, 0, 2039, 0, 15774, 35952, 29633, 32069, 26614, 19840, 11069, 4188, 3144, 4032, 4884, 2755, 7536, 12963, 14266, 24113, 31720, 25324, 33482, 16460, 0, 2820, 0, 1497, 402, 531, 51, 61, 172, 97, 199, 31, 315, 0, 1661, 4313, 3733, 5101, 3256, 6500, 13096, 13002, 22018, 31209, 26641, 35519, 16296, 0, 3183, 37, 1280, 1116, 0, 2080, 0, 16198, 36602, 29902, 33788, 27797, 22784, 14770, 6906, 4797, 4095, 4262, 5458, 1913, 8235, 13749, 20443, 30302, 28602, 29993, 28671, 30368, 27675, 32785, 15608, 0, 3907, 0, 16767, 36236, 29776, 33583, 27639, 22264, 15789, 8883, 4967, 3763, 4097, 5679, 2568, 7356, 13770, 15304, 27553, 27858, 35346, 16309, 0, 2999, 0, 562, 856, 0, 2118, 0, 16381, 36364, 29946, 33246, 29108, 23012, 19956, 20244, 21007, 19038, 23160, 10591, 5318, 15064, 13744, 27279, 28794, 35250, 15994, 0, 3288, 0, 956, 1013, 0, 2431, 0, 16293, 36751, 30546, 33303, 31166, 25890, 22200, 14895, 4211, 4450, 4252, 5628, 2419, 7045, 14023, 14089, 26339, 28598, 34929, 15748, 0, 3076, 0, 1116, 1078, 0, 2695, 0, 16328, 36429, 30074, 32744, 24464, 20943, 14289, 4433, 4458, 4165, 5727, 2287, 7187, 13897, 14948, 27807, 29448, 35820, 16096, 0, 3138, 302, 1950, 331, 1564, 0, 2579, 0, 16027, 36477, 30071, 33566, 26994, 23319, 20089, 10237, 4080, 4226, 4399, 3463, 4767, 2371, 6793, 0, 22315, 20314, 0, 4000, 0, 2217, 582, 1717, 0, 2817, 0, 16404, 36905, 30394, 33981, 30969, 30873, 24963, 16758, 10270, 4218, 4381, 1900, 7401, 18573, 21687, 34819, 15586, 0, 2741, 120, 1834, 1200, 1424, 1467, 1048, 667, 756, 630, 561, 827, 265, 1328, 0, 6002, 11074, 4214, 4652, 4509, 5124, 2534, 8081, 15815, 14979, 27771, 28926, 34930, 17220, 0, 3537, 0, 1384, 1059, 0, 2503, 0, 16379, 36347, 30168, 32247, 23351, 21585, 14651, 5393, 4472, 4910, 5228, 5738, 2213, 9038, 15141, 17253, 22099, 20615, 20949, 21543, 19763, 23733, 10571, 0, 738, 1771, 0, 16124, 35769, 30547, 30147, 23126, 21296, 12232, 5133, 4246, 4568, 5934, 3354, 7790, 14843, 14058, 19895, 25857, 35085, 14972, 0, 3168, 505, 2030, 901, 1957, 0, 2676, 0, 16265, 36431, 29788, 32693, 30687, 31041, 30992, 30607, 31565, 29680, 33472, 21779, 15778, 25356, 35562, 16623, 0, 3428, 330, 2113, 1204, 1920, 1251, 2008, 75, 2708, 0, 16152, 35771, 29300, 32806, 30283, 30748, 24784, 15881, 6548, 1728, 3564, 1780, 6727, 16680, 16292, 31996, 16623, 0, 3257, 0, 1982, 1109, 1738, 1177, 2019, 514, 3318, 0, 16101, 34284, 27819, 27398, 22727, 15631, 4981, 3441, 3465, 4165, 2871, 7368, 14452, 16517, 24683, 33039, 29734, 36772, 16248, 0, 1693, 1659, 0, 16355, 36900, 30245, 32387, 29750, 29819, 29013, 27921, 23691, 21618, 12290, 3158, 3399, 3539, 3877, 3819, 3383, 4541, 2186, 6636, 0, 22412, 20383, 0, 3612, 70, 842, 2018, 0, 15966, 35135, 27987, 31555, 28644, 28150, 25020, 25428, 11248, 0, 3746, 1557, 2941, 0, 6935, 20029, 24129, 31171, 29448, 36006, 16006, 0, 2369, 14, 1654, 1478, 96, 2772, 0, 15362, 34375, 28902, 31031, 30971, 28980, 34205, 15838, 0, 2945, 0, 5048, 16331, 24733, 28990, 29912, 31974, 29412, 36256, 16294, 0, 2933, 0, 2394, 465, 3431, 0, 15918, 36217, 29400, 31128, 28879, 27334, 25291, 9466, 0, 1779, 1095, 635, 11059, 23379, 26350, 29645, 29621, 30690, 30300, 30805, 29908, 31654, 28210, 35258, 14000, 1526, 0, 22156, 16745, 9519, 38367, 26086, 29747, 22054, 9098, 0, 3474, 0, 8898, 21014, 24273, 28528, 29846, 29352, 31444, 28935, 35898, 16249, 0, 2533, 0, 1841, 868, 2232, 871, 2836, 0, 16547, 35490, 27056, 30046, 22272, 18157, 19090, 18827, 18575, 19484, 17349, 24597, 31305, 30456, 31226, 32433, 30028, 36434, 16524, 0, 2076, 0, 478, 2816, 0, 16154, 36292, 30183, 32634, 28146, 30522, 17886, 3259, 4456, 3240, 13825, 22122, 25016, 29858, 30487, 32071, 31596, 33579, 30171, 36702, 16330, 0, 2458, 0, 967, 0, 963, 0, 2289, 0, 16002, 34094, 28667, 19288, 4634, 3891, 6848, 16174, 23886, 29063, 30518, 31508, 31832, 31742, 33305, 29895, 36469, 16276, 0, 2475, 0, 1402, 0, 2795, 0, 16484, 36452, 30499, 33138, 31475, 30800, 27429, 13535, 2631, 9739, 15845, 22940, 28743, 28949, 29449, 28575, 30125, 27330, 32879, 14711, 0, 2485, 0, 1565, 0, 2911, 0, 16675, 36563, 30423, 33436, 31296, 31540, 28193, 12784, 2773, 8696, 14901, 21664, 27249, 30588, 31605, 32000, 31588, 31619, 32421, 32247, 32766, 32174, 33419, 31107, 35756, 18316, 0, 18317, 35418, 30628, 32651, 31806, 31635, 32963, 29985, 36145, 16910, 6369, 23483, 24932, 29928, 30249, 30678, 30501, 30502, 31141, 31830, 31940, 32071, 31675, 31565, 31930, 32240, 32275, 32115, 32088, 31563, 31190, 32102, 31092, 31452, 27302, 20083, 10457, 2015, 9638, 15903, 21414, 28280, 29882, 30980, 31497, 30911, 31115, 32143, 31790, 31970, 31865, 31931, 31871, 32015, 32201, 32140, 31867, 31683, 31584, 32008, 30718, 28946, 19272, 11041, 6219, 5699, 13297, 17381, 23058, 26604, 28413, 29035, 28596, 29814, 30338, 30016, 30299, 30842, 30500, 30335, 30568, 30248, 29969, 30238, 29943, 30442, 30458, 31099, 28800, 27595, 19421, 12678, 14540, 13900, 13730, 14769, 12259, 20958, 30225, 27807, 29711, 29438, 29829, 30268, 30403, 30270, 30073, 29927, 30125, 30359, 30264, 29994, 30213, 30427, 30468, 28715, 29295, 21876, 12744, 8342, 6456, 6418, 13097, 20375, 21643, 26415, 26348, 26959, 27862, 27931, 28212, 28497, 29126, 29152, 29273, 29321, 29294, 29338, 29279, 29364, 29215, 29845, 30420, 25063, 21111, 13674, 6690, 7549, 7096, 8467, 12354, 18858, 24571, 26705, 27194, 27662, 27934, 28249, 28720, 29140, 29134, 29077, 29411, 29628, 29436, 29715, 30283, 30002, 29862, 29227, 29131, 25987, 19376, 15195, 8559, 6580, 7917, 7507, 14879, 18531, 17856, 17764, 18559, 16584, 23502, 30674, 28719, 29827, 29254, 29391, 29384, 29445, 29719, 30219, 30091, 29467, 30683, 27078, 25210, 15718, 7280, 7851, 5594, 8225, 6108, 10343, 14769, 19072, 24756, 25846, 26845, 26982, 28499, 28910, 29212, 29204, 29303, 29276, 29534, 29574, 29667, 30139, 30103, 30352, 29701, 30970, 28605, 33321, 17858, 2871, 9042, 4580, 8483, 17339, 23105, 27385, 28761, 27727, 28296, 28770, 29468, 29895, 29963, 29611, 29618, 29779, 29703, 30044, 30336, 30266, 29745, 30899, 26234, 22061, 14178, 6260, 6387, 5613, 7610, 4089, 8068, 14591, 18613, 26328, 28554, 28127, 28331, 28962, 28784, 28838, 28860, 28735, 29232, 29886, 30094, 30052, 30026, 30203, 30284, 27987, 23279, 22100, 13229, 4856, 6431, 6992, 5291, 9025, 17541, 23129, 28035, 29361, 28543, 28937, 29603, 29843, 29935, 29807, 29790, 29699, 29659, 29715, 30126, 30181, 30575, 29816, 31434, 26147, 23488, 15691, 6047, 7548, 6946, 6643, 7980, 4833, 15897, 29443, 27863, 29047, 29289, 30446, 30314, 30368, 30157, 30263, 30073, 29896, 29929, 30190, 30069, 30427, 30062, 31732, 26307, 24055, 16053, 6005, 6747, 5387, 8458, 4814, 9655, 13980, 17778, 25973, 27779, 28864, 28805, 30113, 30068, 30115, 29992, 29916, 29766, 29794, 29838, 29701, 29993, 29424, 30568, 26729, 21316, 13280, 5679, 5980, 5646, 8077, 4079, 8939, 14081, 17683, 25791, 27172, 28618, 28709, 29788, 29932, 29795, 29654, 29897, 29906, 29920, 29923, 30062, 30500, 30305, 31118, 28745, 25721, 15178, 6459, 6968, 5952, 6382, 7946, 4663, 9098, 15191, 13094, 14490, 13128, 14971, 11697, 22027, 32170, 29352, 30670, 29307, 30131, 29842, 30219, 30769, 30487, 31426, 28656, 26476, 15886, 6471, 6874, 6316, 8267, 6235, 6520, 12518, 14671, 20904, 28693, 28388, 28763, 29472, 30096, 30289, 30200, 30210, 29953, 29922, 30086, 30379, 30499, 30536, 30695, 30636, 30902, 30336, 31392, 29460, 33346, 19697, 1683, 10190, 12970, 17386, 24519, 27543, 28805, 28776, 29889, 29975, 30165, 30180, 30236, 30007, 29837, 30182, 30086, 30045, 30219, 30754, 29757, 27205, 15714, 6127, 6340, 6290, 6142, 8395, 4981, 8840, 13989, 17217, 25730, 27503, 28688, 29033, 30032, 30115, 30122, 30116, 30129, 30088, 30203, 29920, 30435, 29938, 31523, 26160, 23486, 15367, 5035, 7040, 5580, 7051, 6261, 3028, 9620, 15665, 21235, 28481, 28288, 28827, 29616, 30125, 30420, 30297, 30442, 30297, 30262, 30158, 30293, 29836, 30087, 29723, 31016, 25687, 23415, 14973, 5231, 6941, 6314, 7690, 6895, 7724, 6500, 8617, 4456, 18146, 32427, 28971, 31208, 30094, 30602, 30404, 30298, 30271, 30195, 30267, 30021, 30280, 29755, 30152, 25377, 21414, 11969, 4892, 6577, 7538, 3918, 7013, 12728, 16773, 27105, 29268, 29300, 29253, 29897, 30276, 30728, 30415, 30643, 30404, 30339, 30167, 30100, 30171, 30406, 29798, 31000, 28760, 33231, 18322, 2485, 9120, 5457, 8208, 11912, 15953, 25636, 29580, 29378, 29499, 29921, 30451, 30770, 30876, 30694, 30732, 30461, 30601, 30460, 30337, 30055, 29896, 29731, 29498, 28343, 24862, 17557, 8989, 5087, 8430, 4638, 7525, 13262, 16472, 27392, 29485, 29387, 29607, 29480, 29590, 29480, 29610, 29391, 30091, 30910, 30551, 30665, 30291, 29916, 30292, 29540, 29732, 25689, 19753, 10634, 5751, 9632, 4639, 7369, 17437, 22699, 28047, 29820, 29419, 29642, 30044, 30600, 30800, 30811, 31037, 30923, 30727, 30576, 30665, 30757, 30517, 30396, 30622, 30250, 29758, 25769, 23278, 23918, 23702, 23644, 23998, 23132, 26257, 30309, 29739, 30221, 30334, 30474, 30678, 30995, 31108, 30997, 30847, 30787, 30843, 30835, 30574, 30544, 30713, 30727, 30654, 29566, 24264, 16254, 8720, 6484, 8930, 6396, 10131, 17570, 25107, 30745, 29943, 30450, 30189, 30469, 30717, 30788, 30891, 30877, 30922, 30907, 30920, 30914, 30917, 30926, 30852, 30551, 29409, 25182, 13401, 6306, 6741, 8527, 6012, 10259, 14761, 17160, 28038, 30478, 30083, 30083, 12706, 25760, 22450, 11337, 1184, 3837, 0, 470, 1056, 3629, 4108, 3677, 1767, 2568, 1041, 0, 124, 0, 32, 0, 0, 28, 0, 119, 0, 1239, 4028, 5474, 4994, 8193, 9847, 15080, 21082, 19687, 22473, 25434, 26513, 27635, 28270, 28185, 28063, 28414, 27696, 29168, 24377, 20176, 22292, 21689, 21592, 21041, 21427, 21528, 21735, 22306, 21944, 20645, 22078, 22790, 23416, 23915, 25743, 22984, 18562, 18503, 19652, 20407, 18202, 19336, 20896, 21055, 22585, 24418, 22613, 23110, 25211, 26834, 28088, 25413, 26012, 13365, 5372, 7934, 5554, 6688, 5996, 6527, 5939, 6903, 4029, 2120, 3784, 3068, 2583, 1739, 1351, 1257, 1546, 1933, 1838, 466, 0, 39, 0, 12, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 80, 0, 322, 0, 5770, 15008, 18373, 22770, 24071, 24417, 25685, 25131, 25320, 25941, 26901, 27885, 29350, 29243, 25481, 23464, 20523, 17285, 20750, 20687, 24541, 14290, 9120, 19768, 21694, 23758, 23238, 22996, 24029, 21854, 26320, 11631, 0, 1381, 0, 638, 82, 75, 843, 2033, 2818, 3698, 3501, 3584, 3388, 3288, 3017, 2961, 3134, 3416, 2939, 2501, 2390, 2144, 3006, 3797, 4020, 5544, 3482, 9974, 18952, 18564, 21149, 24689, 22520, 29133, 13004, 0, 1616, 0, 467, 0, 95, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 121, 0, 433, 0, 3693, 9499, 9360, 8580, 9391, 11643, 11597, 11058, 15944, 19841, 18454, 17904, 17910, 18368, 19392, 19852, 19394, 18750, 17682, 18224, 18433, 17869, 18665, 19661, 19379, 19471, 19511, 19324, 19775, 18268, 17089, 17473, 17536, 16655, 17733, 13954, 9518, 11669, 9658, 10127, 12060, 10516, 4050, 0, 4594, 12644, 16987, 18464, 12559, 14011, 6401, 0, 820, 0, 239, 0, 63, 0, 217, 775, 409, 0, 340, 195, 0, 24, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 272, 0, 946, 0, 8598, 20006, 17531, 17319, 15457, 16386, 15945, 16118, 15313, 17670, 18526, 20617, 8822, 0, 2402, 3030, 6627, 6736, 5121, 4914, 3747, 3661, 2580, 1747, 707, 0, 89, 0, 24, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 44, 72, 1530, 1056, 1751, 4995, 5630, 7048, 7204, 8664, 3723, 0, 459, 0, 131, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 83, 0, 411, 0, 1436, 0, 11763, 27725, 23827, 24632, 22985, 25439, 25492, 24884, 24997, 24610, 25183, 24471, 25063, 26255, 24584, 23622, 23676, 22171, 21285, 21429, 20739, 20445, 19876, 19992, 19217, 18585, 18476, 19284, 18932, 22269, 21989, 18551, 20410, 18452, 16463, 15888, 15802, 15835, 15767, 15600, 16086, 15073, 16995, 13312, 22857, 15282, 0, 5774, 1619, 329, 699, 1891, 2189, 2220, 2247, 2484, 1608, 115, 15, 0, 0, 64, 404, 2393, 1357, 0, 179, 0, 52, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 104, 0, 408, 0, 2266, 756, 4064, 15633, 19072, 21770, 23306, 23948, 25197, 23736, 24497, 19165, 17877, 8396, 0, 1078, 0, 243, 0, 0, 315, 0, 3308, 9272, 3135, 0, 310, 0, 100, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 31, 159, 78, 0, 9, 0, 2, 0, 0, 5, 0, 24, 0, 81, 0, 1093, 4835, 6288, 5671, 6522, 5040, 7721, 2537, 17582, 20260, 7282, 8608, 463, 238, 0, 38, 0, 0, 5, 0, 0, 0, 0, 8, 0, 37, 0, 131, 0, 1179, 3575, 3120, 2763, 1554, 1970, 0, 9636, 24907, 26188, 28631, 28234, 29488, 28763, 28265, 27608, 26023, 25182, 25445, 25242, 25487, 25110, 25822, 23438, 20356, 20285, 19013, 18508, 17723, 17119, 16697, 16310, 16172, 16317, 17274, 18919, 19721, 19493, 16599, 15596, 19244, 10929, 5003, 7502, 6661, 6884, 6151, 6518, 17073, 24275, 24976, 26917, 25159, 19450, 8997, 3489, 2710, 1876, 1847, 2051, 1883, 1913, 1911, 1882, 1964, 1805, 2128, 1006, 0, 460, 276, 0, 34, 0, 11, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 23, 0, 192, 827, 1816, 3018, 1633, 7428, 13717, 15847, 21007, 23296, 23642, 21416, 18785, 17089, 16302, 16805, 16311, 18349, 21186, 22552, 19730, 17013, 6386, 0, 7364, 10793, 8836, 9272, 3936, 0, 477, 0, 140, 0, 27, 0, 1, 0, 11, 0, 38, 0, 663, 1858, 2748, 3529, 3258, 3311, 3504, 3654, 3781, 3685, 3716, 3596, 2509, 1894, 1894, 1622, 1710, 1459, 3097, 3932, 4586, 4000, 5870, 2406, 12308, 25906, 22046, 20879, 24687, 9918, 0, 1158, 0, 333, 0, 70, 0, 0, 0, 0, 0, 0, 6, 0, 34, 0, 95, 0, 801, 2480, 1630, 2344, 0, 10313, 24274, 22415, 25447, 25274, 25875, 25584, 25836, 26001, 26315, 26352, 25941, 23789, 22601, 23308, 23246, 22388, 23962, 24632, 23864, 21914, 19688, 19157, 18161, 18040, 17932, 17761, 17395, 17697, 17203, 18096, 16467, 19671, 9693, 3259, 9134, 6090, 6320, 6280, 6428, 7092, 4967, 797, 286, 978, 2665, 2316, 1371, 1334, 849, 1214, 1711, 2047, 1812, 1522, 1960, 1966, 543, 0, 55, 0, 48, 0, 249, 794, 2421, 1300, 0, 170, 0, 49, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 37, 0, 199, 0, 1132, 0, 8007, 21233, 20528, 21420, 20828, 21280, 20791, 21596, 19051, 16155, 16279, 17283, 19917, 20953, 19122, 14418, 4529, 0, 3401, 14441, 18790, 19527, 15266, 5657, 1486, 0, 173, 0, 34, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 7, 0, 24, 0, 199, 448, 376, 405, 401, 382, 439, 215, 0, 199, 597, 228, 0, 0, 46, 0, 1074, 6234, 9094, 11926, 5185, 0, 746, 0, 195, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 32, 0, 164, 0, 544, 902, 2893, 4474, 3434, 4252, 3175, 4928, 1573, 12420, 23200, 20199, 22071, 22143, 23468, 22500, 20877, 22843, 24062, 23848, 24893, 23465, 24606, 23903, 21178, 19759, 18515, 17722, 16665, 16127, 15745, 15270, 16044, 16557, 16165, 17545, 16395, 17665, 11099, 5187, 8005, 7319, 8672, 8814, 5604, 998, 8824, 19159, 20356, 20006, 20787, 19197, 22455, 11869, 1861, 3608, 752, 1934, 1596, 863, 0, 107, 0, 59, 0, 119, 0, 833, 1360, 374, 192, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 57, 0, 160, 0, 1489, 4606, 3229, 5763, 1114, 7363, 20646, 20971, 23350, 9157, 0, 1933, 570, 1146, 921, 562, 139, 283, 489, 0, 2158, 5030, 2547, 1505, 1683, 1663, 1568, 1845, 831, 0, 102, 0, 29, 0, 5, 0, 0, 0, 0, 3, 0, 16, 0, 56, 0, 411, 692, 456, 908, 813, 458, 1095, 2447, 2710, 2968, 2641, 273, 3626, 8560, 9227, 9698, 12313, 13191, 12198, 12959, 12630, 12460, 12512, 12458, 12527, 12421, 12669, 11071, 3939, 0, 167, 0, 52, 0, 9, 0, 0, 0, 0, 49, 0, 240, 0, 837, 0, 7514, 21314, 22800, 27236, 30362, 31025, 30856, 31346, 31548, 31996, 32326, 31497, 30171, 27492, 26478, 26711, 26255, 26145, 25988, 25563, 25156, 25289, 25209, 25282, 25186, 25352, 24856, 24417, 24103, 23459, 23556, 23576, 24104, 24602, 24859, 25195, 24324, 21504, 19504, 19278, 18965, 19941, 21304, 22936, 24458, 22768, 21090, 25117, 24495, 20115, 8238, 1880, 2901, 1700, 3811, 3316, 5347, 6432, 5307, 1991, 0, 2599, 5738, 4915, 4984, 4934, 4865, 5091, 4628, 5575, 2465, 0, 306, 0, 87, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 75, 0, 250, 0, 3405, 15416, 19812, 18479, 18276, 16906, 17858, 16008, 19197, 6583, 3940, 19007, 19603, 22552, 24287, 23623, 24074, 26098, 24988, 22972, 21396, 20245, 20491, 23346, 22809, 22777, 24493, 21205, 20225, 19206, 21272, 14104, 6808, 6681, 3291, 3668, 3274, 3329, 3139, 3225, 3145, 3274, 3046, 3498, 2015, 588, 1524, 1933, 2092, 2063, 2195, 2211, 1688, 319, 3336, 8024, 11633, 13358, 14588, 22114, 26490, 24246, 24221, 26684, 28858, 29336, 29366, 29962, 30072, 30298, 31517, 31031, 29823, 26758, 25187, 19917, 20221, 9041, 0, 1138, 0, 320, 0, 62, 0, 0, 0, 11, 0, 58, 0, 198, 0, 3011, 12765, 18548, 21312, 22266, 21350, 22577, 24929, 26370, 26664, 25876, 26269, 22384, 18865, 19347, 18553, 18221, 17970, 18215, 17875, 17427, 16893, 16614, 16941, 16317, 15817, 15334, 16180, 17344, 17573, 18236, 18734, 19100, 18861, 19074, 18760, 19294, 18336, 20274, 13308, 2183, 1395, 1437, 1855, 2301, 2342, 2620, 3133, 1819, 1188, 503, 0, 410, 2658, 2452, 1302, 2280, 1800, 1111, 994, 925, 199, 0, 0, 73, 0, 345, 363, 0, 55, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 25, 0, 55, 72, 2588, 5672, 5741, 7420, 4884, 10728, 22248, 22524, 22363, 22738, 22643, 22640, 22748, 22490, 23042, 21062, 18839, 21515, 20223, 20401, 20195, 15665, 17301, 7784, 2840, 9833, 10357, 12818, 11056, 12311, 5887, 0, 644, 0, 182, 0, 34, 0, 0, 0, 11, 0, 44, 0, 172, 0, 2185, 6407, 5514, 2925, 7813, 9500, 9555, 11841, 11054, 11358, 11394, 11004, 11949, 9048, 8127, 9047, 7013, 5500, 1792, 354, 619, 2048, 2673, 5575, 3825, 0, 193, 0, 60, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 74, 0, 242, 153, 8578, 16048, 18496, 21083, 20183, 20669, 20359, 20622, 20264, 21340, 22799, 23198, 23571, 23368, 22950, 22120, 21897, 21131, 20401, 20723, 20691, 20924, 20235, 19747, 19749, 18777, 18349, 18122, 18222, 18674, 18256, 17688, 18130, 17823, 17199, 15342, 10460, 9480, 9746, 11224, 9032, 10197, 12120, 14185, 20127, 20529, 19352, 17813, 18467, 17842, 18729, 17232, 20143, 10564, 454, 3250, 406, 34, 0, 0, 6, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 40, 0, 197, 0, 896, 0, 3795, 9951, 14660, 20107, 15163, 4134, 0, 392, 0, 107, 0, 15, 0, 0, 29, 159, 2590, 4954, 4758, 3664, 3498, 1443, 0, 200, 0, 76, 7, 24, 0, 1, 0, 0, 0, 0, 7, 0, 37, 0, 130, 0, 1042, 2300, 1890, 2173, 2044, 2055, 2017, 2021, 2024, 1856, 1708, 1649, 1613, 1594, 1518, 1441, 1422, 1616, 1867, 2036, 1980, 2709, 5909, 9766, 8580, 8233, 9745, 8992, 9736, 8698, 10562, 4653, 0, 579, 0, 165, 0, 34, 0, 8, 0, 29, 0, 312, 1440, 2480, 2408, 1915, 12020, 20091, 23416, 26920, 25331, 25400, 25123, 22176, 19820, 19620, 19568, 19873, 19966, 19855, 19256, 19084, 18755, 18846, 18930, 18688, 18844, 18836, 18792, 18783, 18831, 18721, 18958, 18220, 17573, 17246, 18981, 19915, 17938, 18254, 16986, 16460, 14720, 13020, 13509, 10811, 13739, 15606, 18752, 18477, 22712, 24000, 22737, 11616, 882, 2915, 0, 1746, 2144, 1749, 2008, 1718, 2001, 1215, 29, 35, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 190, 0, 661, 0, 6181, 18853, 21117, 22483, 22730, 22882, 22924, 23283, 23176, 23722, 23797, 22857, 24818, 24070, 23749, 9720, 0, 7637, 17860, 14018, 13379, 14329, 7309, 1940, 0, 207, 0, 44, 0, 23, 0, 80, 0, 277, 0, 2409, 6270, 5153, 4892, 4930, 4831, 5041, 4654, 5419, 2825, 0, 1287, 1467, 1763, 754, 0, 7, 431, 3267, 8962, 9716, 8485, 6592, 9088, 13302, 12149, 14843, 19559, 21608, 27597, 18337, 11698, 6660, 0, 962, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 57, 0, 283, 0, 992, 0, 7926, 17663, 14838, 17510, 16855, 17928, 18571, 18876, 19270, 19431, 19789, 19997, 20166, 20291, 20375, 20737, 20656, 21557, 23856, 24150, 23558, 24031, 23311, 23260, 20214, 25491, 27988, 24004, 13697, 5448, 6853, 5995, 6182, 5308, 6004, 5683, 2107, 0, 240, 0, 67, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 38, 0, 40, 297, 5618, 14010, 7282, 15321, 28184, 26516, 21257, 15779, 17541, 16987, 16547, 16181, 16147, 16768, 17794, 18133, 18624, 18736, 19253, 19641, 20221, 20471, 20382, 20494, 20279, 20709, 19871, 21711, 20055, 26761, 26382, 19699, 22117, 21631, 19063, 17894, 11696, 4483, 4112, 2428, 1303, 0, 172, 0, 38, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 31, 0, 153, 0, 536, 0, 4394, 9580, 8452, 8278, 9677, 6225, 18398, 30875, 22218, 21584, 21178, 20698, 20600, 20220, 20614, 20612, 20152, 20205, 20340, 20638, 20965, 23174, 30120, 31980, 32144, 29172, 37029, 15571, 0, 0, 15421, 34008, 22774, 19129, 18505, 23229, 21126, 17480, 5680, 126, 750, 0, 161, 0, 36, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 129, 0, 430, 0, 3843, 10014, 7531, 9730, 13605, 18111, 26761, 30427, 28717, 28671, 24946, 22351, 22571, 21472, 21914, 22043, 21905, 21344, 20938, 21436, 21589, 21369, 21415, 21180, 21467, 21234, 21479, 21978, 21808, 21908, 21831, 21933, 21765, 21959, 19996, 19793, 19926, 19190, 8456, 0, 4131, 4590, 4994, 2042, 0, 254, 0, 75, 0, 14, 0, 0, 0, 1, 0, 10, 0, 36, 0, 240, 240, 0, 36, 0, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 102, 0, 296, 0, 2906, 7102, 0, 9920, 27324, 29531, 31529, 30956, 31280, 31179, 31067, 31473, 30588, 32262, 29169, 35913, 16146, 0, 2256, 0, 1134, 1895, 3955, 3297, 3599, 2790, 3306, 1443, 3852, 0, 16782, 35073, 27818, 28655, 22054, 22364, 23653, 20001, 6623, 0, 694, 0, 181, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 105, 0, 322, 0, 3190, 9288, 4798, 9627, 15717, 19710, 27828, 30558, 31347, 30268, 29207, 26402, 23155, 21905, 22075, 21798, 21648, 22142, 23624, 24235, 24683, 23374, 25229, 22271, 33305, 17536, 0, 3403, 0, 2017, 1674, 2870, 2642, 1528, 1952, 1713, 1873, 1731, 1923, 1299, 403, 945, 0, 2277, 6850, 7775, 8167, 8302, 8872, 8795, 9020, 7474, 5598, 6675, 7405, 8214, 8700, 8169, 7417, 6650, 4750, 4999, 4915, 5909, 2870, 0, 371, 0, 104, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 163, 0, 539, 0, 4521, 10074, 4279, 8760, 14710, 19107, 25721, 30318, 30763, 26748, 25738, 21891, 18895, 19521, 19405, 19231, 19891, 18431, 21248, 15829, 29745, 18033, 0, 4696, 1512, 5281, 5162, 5092, 5775, 5829, 5917, 6127, 6151, 4856, 5184, 0, 13582, 25385, 14090, 6237, 768, 1909, 614, 903, 705, 797, 289, 0, 35, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 109, 0, 499, 0, 1983, 0, 11685, 28965, 24325, 26037, 21332, 19025, 19221, 18614, 19794, 20208, 20578, 20922, 21017, 20962, 21243, 21572, 21837, 21775, 21766, 21643, 20775, 21489, 22471, 22644, 27742, 20929, 34660, 12422, 12324, 35423, 21062, 26689, 24301, 24890, 24598, 21924, 19470, 20332, 19622, 20510, 19124, 21738, 13097, 3631, 7350, 2351, 0, 234, 0, 151, 0, 281, 0, 2094, 4791, 3842, 4251, 3958, 4475, 1704, 0, 200, 0, 57, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 103, 0, 292, 0, 3353, 11141, 4450, 8221, 16035, 15380, 18539, 18860, 19187, 19496, 19709, 19862, 20750, 20796, 21076, 21245, 21451, 21585, 21634, 21452, 21837, 21039, 23612, 25825, 24829, 23142, 21351, 21020, 19519, 20697, 21754, 20199, 11196, 6109, 6861, 5544, 5759, 5151, 6622, 8720, 6012, 4220, 5010, 4119, 4802, 1911, 0, 227, 0, 67, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 438, 0, 1506, 0, 12442, 28816, 19438, 18068, 18009, 18403, 17932, 18290, 19011, 19838, 20618, 20808, 21025, 20779, 21036, 21187, 21365, 20914, 22899, 26560, 25798, 26292, 24456, 27335, 27085, 33345, 19627, 0, 18629, 34932, 25448, 19740, 15924, 17806, 19243, 11335, 6692, 4341, 0, 217, 0, 60, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 147, 0, 493, 0, 4172, 9760, 4641, 2635, 2205, 531, 0, 32, 0, 8, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 79, 0, 267, 0, 2188, 4775, 2083, 1288, 1314, 680, 48, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 88, 0, 288, 0, 2339, 4261, 0, 6204, 15984, 17457, 17287, 17438, 17222, 17538, 16817, 21753, 37370, 15500, 0, 3032, 227, 2605, 2112, 2471, 2234, 2285, 2782, 3209, 3137, 3373, 4195, 4500, 4193, 4592, 1714, 4734, 0, 15678, 32807, 22287, 25785, 25236, 22486, 22596, 8420, 788, 0, 10070, 9920, 0, 5958, 0, 352, 0, 66, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 127, 0, 457, 0, 4165, 9244, 10541, 12850, 10239, 9002, 2931, 6198, 22911, 21972, 16411, 18675, 17980, 17749, 17582, 18728, 19000, 19810, 21235, 21977, 23687, 23396, 22909, 24555, 23688, 21992, 22438, 23736, 24820, 29860, 28939, 35673, 16179, 0, 2304, 0, 531, 1089, 0, 6444, 6629, 0, 1529, 65, 828, 444, 472, 223, 218, 260, 85, 0, 8, 0, 1, 2, 0, 22, 0, 81, 0, 530, 530, 0, 81, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 83, 0, 276, 0, 2607, 7336, 6724, 3625, 1670, 0, 13414, 21429, 17289, 19638, 18543, 19581, 19646, 19638, 19721, 19545, 19851, 19257, 21151, 22935, 22545, 22724, 22267, 22279, 21851, 24628, 27149, 24741, 27539, 32784, 30795, 23864, 22747, 13765, 5815, 7810, 5115, 6200, 5928, 6160, 2958, 0, 277, 0, 78, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 162, 0, 653, 0, 6489, 7136, 3492, 0, 14317, 29687, 24169, 23405, 18579, 20479, 19563, 21278, 23313, 25140, 27063, 27712, 27739, 27366, 27637, 26181, 23214, 21469, 20811, 20268, 22361, 24614, 26612, 23505, 31017, 19087, 0, 18996, 33936, 23628, 24946, 14906, 6953, 9348, 7958, 9059, 7871, 9686, 4243, 0, 529, 0, 151, 0, 30, 0, 0, 0, 0, 3, 0, 12, 0, 38, 0, 444, 1526, 616, 0, 69, 0, 21, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 42, 0, 105, 661, 8227, 8417, 3423, 2430, 0, 2125, 11597, 17440, 17668, 18298, 18003, 19807, 20255, 23072, 23261, 21401, 22177, 21800, 21984, 21916, 21962, 21769, 21819, 23652, 27961, 23301, 32044, 19235, 0, 19399, 33264, 26662, 26473, 24415, 26163, 23739, 19952, 9656, 3727, 6890, 2106, 0, 186, 0, 62, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 74, 0, 366, 0, 1288, 0, 10855, 27395, 25502, 22392, 18647, 20257, 19499, 19698, 19738, 20149, 20267, 20757, 21228, 21111, 21448, 21142, 21293, 21741, 21555, 21152, 20639, 20904, 20554, 22597, 26510, 24103, 26374, 30477, 21988, 21456, 14053, 5777, 8255, 6389, 6815, 5964, 5753, 5788, 4489, 3731, 3848, 3938, 3629, 4335, 1928, 0, 238, 0, 68, 0, 11, 0, 0, 27, 0, 100, 0, 818, 1996, 2033, 842, 0, 103, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 162, 0, 582, 0, 4201, 6600, 1948, 305, 2941, 15104, 19036, 18343, 19022, 18635, 18152, 18538, 20156, 20832, 20935, 21126, 21506, 21546, 21422, 21386, 21518, 21702, 21819, 21683, 21942, 21472, 22320, 20634, 26292, 30323, 16367, 5516, 3336, 2875, 2824, 2606, 2312, 1969, 2116, 901, 0, 110, 0, 31, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 191, 0, 667, 0, 4893, 8080, 2404, 3002, 2282, 2983, 2057, 3572, 637, 10225, 19934, 17539, 20708, 21182, 20868, 20122, 20574, 21052, 21258, 21013, 21211, 21377, 21364, 21212, 21419, 21482, 27775, 21545, 34290, 13887, 10549, 31533, 6951, 3962, 4052, 6030, 14176, 19437, 10748, 5811, 7821, 5111, 7521, 3920, 0, 519, 0, 151, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 11630, 8074, 19192, 29488, 25144, 26928, 23844, 25560, 9572, 0, 932, 0, 0, 2918, 8724, 7436, 8324, 7992, 8530, 10130, 9630, 9660, 9624, 9534, 10326, 10318, 10378, 9896, 10700, 9538, 12560, 4490, 3016, 12614, 11238, 12566, 11578, 11718, 11632, 11866, 12104, 12070, 12000, 12190, 11806, 12596, 9890, 6892, 8846, 9072, 8208, 10218, 12550, 12362, 11748, 11698, 11846, 12224, 12110, 10914, 11758, 8420, 14882, 2768, 11280, 27998, 22324, 32052, 27504, 26262, 24958, 19828, 25290, 26892, 24638, 24486, 22016, 21898, 28158, 30710, 31742, 28730, 25610, 28498, 27992, 28402, 28108, 28388, 27996, 28724, 26352, 24106, 24488, 23482, 24052, 28258, 24098, 26572, 29444, 22292, 31272, 28730, 19626, 26606, 26020, 17760, 15174, 14088, 8060, 15198, 17732, 17432, 22274, 21850, 19862, 22770, 21076, 32880, 16076, 1532, 14598, 9820, 13350, 12298, 14186, 14412, 14906, 14712, 14528, 14670, 14428, 14842, 14122, 15456, 11468, 9844, 16616, 10584, 24430, 30042, 35884, 26098, 9482, 18552, 16230, 17930, 17594, 18792, 19282, 17678, 17194, 16518, 16030, 16244, 17108, 18822, 18108, 19064, 16608, 17562, 17962, 15088, 15620, 16198, 12582, 9124, 10644, 14972, 14612, 17118, 10192, 21008, 35820, 31288, 33220, 32842, 31764, 34972, 24070, 13932, 9358, 18080, 32684, 31646, 34322, 27792, 33180, 35566, 37352, 39148, 44100, 30170, 20016, 17308, 31296, 32964, 14226, 20696, 16896, 15098, 25094, 35480, 28964, 33836, 29384, 17772, 27020, 34704, 32170, 24368, 14050, 21166, 30774, 28998, 33536, 34590, 32896, 33656, 33008, 33800, 32596, 34836, 27392, 18878, 21770, 17180, 14442, 14938, 14304, 14096, 13650, 12676, 12228, 10600, 9786, 10932, 9814, 10790, 13734, 14724, 17958, 18940, 14580, 16718, 22260, 23382, 23438, 25594, 20396, 16250, 17378, 16716, 16888, 16000, 16282, 15796, 15668, 15898, 15430, 15606, 15848, 15726, 15872, 15636, 16120, 14156, 10332, 12200, 16180, 10200, 8802, 14296, 19192, 20592, 24558, 23222, 34742, 44016, 42606, 30766, 17098, 20958, 18290, 21822, 8578, 0, 2158, 0, 11028, 30066, 29810, 35230, 23606, 16508, 22546, 21470, 22538, 23858, 22630, 24950, 21632, 34506, 43074, 37144, 41130, 39090, 40484, 39164, 41070, 35626, 30984, 30850, 30740, 34678, 35528, 36254, 37272, 38170, 36320, 38030, 34640, 39118, 18318, 0, 13118, 22864, 21872, 23674, 23552, 24276, 24998, 24178, 23726, 18074, 17234, 22192, 20598, 20246, 21114, 19402, 22976, 26106, 26332, 27806, 25982, 24518, 25780, 24022, 22006, 22676, 22234, 22664, 22048, 23682, 24344, 23218, 22598, 22622, 23752, 24070, 24764, 25064, 24980, 25626, 26232, 25730, 25866, 26062, 23832, 22260, 22266, 40554, 33178, 29178, 37426, 41922, 40066, 26434, 35918, 18412, 9630, 20674, 14758, 25286, 15000, 8452, 28644, 28362, 32680, 24668, 24196, 32796, 31100, 32062, 31838, 31296, 32890, 28890, 31420, 18946, 23176, 29792, 29128, 35828, 22092, 32920, 22280, 19810, 40820, 27268, 14888, 19934, 20694, 14374, 11252, 1040, 19380, 25418, 23034, 30114, 17770, 21134, 15536, 27834, 36238, 43188, 25918, 14130, 28446, 24156, 27140, 26144, 27158, 27312, 27316, 27190, 27138, 27274, 27050, 27418, 26626, 30974, 43514, 34346, 35782, 46210, 36152, 22986, 24484, 37156, 37878, 44792, 33520, 21796, 28254, 27934, 28806, 26220, 21522, 24578, 28010, 28612, 29106, 28388, 27380, 24888, 21754, 19572, 19812, 17594, 24360, 39302, 34866, 23314, 26214, 35354, 32448, 23270, 19498, 17866, 18432, 18012, 18484, 17776, 19166, 13808, 4034, 10420, 24682, 29954, 28790, 31572, 24102, 13872, 23982, 38178, 36050, 38918, 45238, 36620, 45800, 35432, 30192, 33018, 31302, 30580, 23898, 13394, 15216, 23768, 26168, 37348, 30526, 29494, 17756, 14326, 23874, 27934, 28256, 29030, 21360, 22284, 34462, 34512, 35192, 34682, 35124, 34584, 35556, 31880, 25264, 27602, 25426, 24940, 22426, 17250, 17940, 14956, 18716, 21998, 21476, 20238, 11278, 7452, 8654, 9174, 8730, 16634, 19194, 14432, 22950, 28190, 27760, 31562, 24374, 17494, 19558, 18532, 18578, 17968, 18108, 17564, 17890, 17384, 18990, 20098, 18340, 18096, 18148, 17992, 18326, 17696, 18916, 15294, 14266, 18030, 16514, 18716, 20308, 20992, 29350, 23918, 33384, 45466, 38622, 40314, 41088, 38184, 38902, 27716, 9706, 0, 19990, 14870, 7266, 39058, 30496, 45048, 20628, 9518, 27750, 25580, 29048, 29210, 27092, 27376, 26504, 35246, 46128, 41836, 44872, 46484, 46238, 46166, 46556, 45668, 47604, 40436, 29504, 32444, 36522, 36822, 35746, 37868, 40554, 42812, 44086, 38868, 45890, 21390, 0, 13606, 26194, 26522, 28214, 28364, 29464, 29274, 30496, 28698, 28474, 23302, 21350, 26810, 25588, 25938, 23230, 27192, 48484, 24194, 15260, 32342, 26072, 30012, 28224, 28490, 28230, 28474, 28032, 28930, 27230, 30264, 18042, 15190, 27592, 27372, 29536, 29556, 30328, 30468, 30952, 31514, 31340, 32168, 29184, 35280, 44984, 44926, 42114, 39426, 41440, 41080, 34606, 34112, 37498, 35000, 33616, 31568, 34604, 28124, 19092, 19562, 16696, 18804, 26398, 32114, 37154, 26716, 23952, 30660, 28114, 29602, 28504, 29588, 28024, 32452, 34372, 24314, 26070, 24246, 37048, 34688, 35744, 33426, 31216, 27180, 11558, 18996, 25154, 16102, 13220, 19918, 19832, 11596, 13594, 23302, 17818, 20946, 20720, 19930, 24990, 34120, 33606, 43356, 30268, 20738, 30264, 28356, 30744, 30456, 31634, 30050, 29802, 31158, 30600, 31052, 30440, 31518, 29492, 33966, 29022, 37098, 36358, 31902, 43508, 21980, 23852, 33436, 30310, 35362, 38916, 49030, 36592, 24750, 30060, 30116, 32682, 29518, 27292, 28326, 29934, 31264, 30034, 28854, 23854, 24518, 19896, 28278, 43422, 33588, 25030, 27506, 25776, 24582, 35082, 38384, 39028, 40638, 40306, 40028, 41022, 38910, 43300, 28778, 13594, 17622, 24370, 34644, 33462, 35974, 28512, 17852, 31400, 33248, 37024, 45472, 44892, 44942, 44444, 25660, 27090, 48668, 25178, 29360, 31288, 29884, 34450, 35782, 30102, 32630, 30878, 23892, 33160, 23482, 18474, 15902, 18114, 18398, 18806, 20378, 30534, 35768, 34456, 34992, 34888, 34588, 35502, 32136, 28008, 27558, 27804, 25838, 25080, 25460, 28084, 21014, 17318, 23414, 23016, 25674, 25350, 23424, 22666, 21368, 24406, 17994, 26244, 9614, 25418, 38608, 20214, 31688, 30008, 27362, 20190, 23090, 24340, 24296, 21902, 20530, 20474, 20242, 21070, 24544, 27726, 28304, 28256, 28250, 28264, 28198, 28496, 26212, 18048, 17682, 19334, 0, 21600, 43684, 37268, 46736, 43836, 46790, 45028, 40512, 35608, 36316, 36140, 34922, 35658, 33890, 33416, 31576, 30554, 23394, 30470, 36038, 46954, 19110, 3216, 28106, 24568, 30352, 23594, 23678, 15052, 34902, 51396, 36942, 42826, 43762, 44252, 43372, 45016, 41864, 48170, 29460, 22016, 24108, 21412, 35244, 34544, 37944, 36736, 40378, 44768, 46528, 38710, 50340, 20070, 2478, 26306, 24672, 28896, 28398, 30218, 30090, 30768, 29558, 29136, 30022, 29746, 27950, 28066, 27482, 28400, 24028, 36108, 49294, 47270, 48044, 52444, 39576, 21840, 22584, 21434, 22290, 21436, 22618, 20554, 25754, 22626, 20656, 28024, 27964, 30184, 30022, 30552, 30840, 31442, 32066, 32706, 30438, 32054, 25802, 36210, 48444, 46160, 48620, 45972, 43924, 34012, 28318, 36644, 30812, 19166, 17886, 19288, 20622, 18670, 16318, 12446, 16858, 17278, 27296, 24372, 24228, 37502, 36198, 36904, 37428, 35370, 39920, 27740, 31280, 26706, 23530, 35540, 21520, 30254, 26092, 34542, 37542, 20416, 31842, 23970, 26274, 31916, 19392, 18808, 13592, 19138, 21794, 16810, 18036, 20614, 19990, 22536, 18176, 29332, 32596, 42454, 23490, 10680, 32104, 25426, 30026, 30576, 31888, 31930, 31716, 31672, 31390, 31518, 31390, 31582, 31324, 31196, 28064, 37212, 49208, 35160, 31098, 28000, 15928, 28780, 36528, 33052, 30526, 37328, 49032, 34644, 26090, 31012, 31838, 30942, 29918, 31288, 31106, 31918, 31762, 30110, 29380, 29426, 23382, 33514, 45040, 39598, 39280, 32260, 27832, 30040, 30896, 27792, 27284, 36974, 40408, 39216, 40566, 38462, 42408, 29604, 16364, 21670, 17812, 27914, 38360, 28714, 21596, 20828, 20002, 21790, 34292, 40114, 42374, 43662, 37566, 33996, 39734, 34910, 22080, 32114, 30910, 17520, 25004, 25368, 21208, 25154, 18436, 17184, 17578, 21452, 15544, 14658, 20936, 19090, 20456, 19316, 19426, 19112, 18820, 19118, 18636, 19476, 17820, 23482, 30568, 29018, 29718, 28758, 26136, 27970, 24472, 23572, 22458, 21248, 24006, 27048, 20574, 20250, 24530, 23102, 18316, 2378, 15010, 24008, 22774, 26408, 26764, 30344, 31450, 28010, 23076, 22216, 22112, 21534, 20054, 20554, 20390, 21738, 21406, 23802, 26828, 25852, 26366, 26016, 26366, 25844, 26812, 24226, 22706, 16958, 28564, 42328, 34740, 34660, 42838, 40120, 40360, 39772, 27672, 32024, 38208, 27480, 25532, 35258, 36606, 35082, 32622, 29488, 32818, 36676, 39232, 38856, 45916, 23606, 12810, 27582, 25932, 25054, 34564, 50082, 47156, 47884, 37104, 36956, 44568, 42426, 43878, 42604, 44136, 41754, 46274, 31398, 15374, 20732, 19124, 28940, 37900, 37938, 37972, 41704, 46780, 40478, 48952, 21410, 0, 15964, 22698, 26812, 26880, 28512, 29076, 29262, 28890, 28074, 28168, 28810, 28186, 27584, 26294, 25460, 20312, 34996, 48092, 46692, 48018, 52662, 35758, 23264, 17826, 6298, 10322, 8200, 9468, 8536, 9500, 8548, 18336, 27612, 27902, 29434, 29544, 30130, 29556, 29670, 31232, 28690, 27514, 32808, 21564, 33556, 43028, 42630, 43134, 30908, 43916, 39680, 29734, 29020, 14866, 27784, 28568, 17354, 32942, 29076, 19334, 13740, 16002, 19996, 23638, 30672, 24408, 30414, 36398, 33366, 34866, 33750, 34968, 33130, 36480, 27596, 26858, 20750, 26438, 38376, 22254, 28408, 27966, 19790, 20224, 23562, 22778, 21044, 33782, 28072, 17114, 21148, 14504, 14282, 17882, 17804, 20976, 22062, 21574, 24000, 31734, 35042, 46346, 22250, 12136, 27848, 24590, 30538, 29524, 31540, 30216, 30506, 28552, 26154, 26800, 26676, 26410, 27122, 25510, 32306, 45816, 36406, 31296, 27828, 28056, 32464, 32752, 35622, 32134, 37122, 41210, 49134, 37316, 24752, 28916, 29682, 31194, 30558, 32070, 32140, 30452, 29040, 27674, 28986, 27648, 39676, 36338, 23872, 28486, 25628, 22288, 20870, 23826, 20710, 21680, 25280, 22826, 21980, 22248, 21848, 22578, 21246, 23834, 16152, 13388, 18888, 18036, 20406, 20928, 20940, 18498, 16698, 22328, 32960, 37734, 41576, 37682, 42504, 29464, 30460, 36506, 29866, 40632, 32904, 10046, 15002, 12716, 7500, 21098, 22546, 20334, 9156, 16494, 11604, 7906, 16206, 16984, 17580, 18272, 15724, 25298, 34610, 31842, 33150, 32558, 32664, 33086, 30486, 23866, 23668, 21564, 18508, 19358, 17502, 15856, 13998, 17174, 23020, 22908, 22124, 14526, 7028, 18122, 18864, 22126, 13156, 9756, 24422, 22886, 26258, 27964, 31754, 26296, 19660, 22102, 21258, 19616, 19404, 19362, 19422, 19212, 20308, 19226, 22438, 22790, 19620, 20668, 20332, 20072, 21072, 18954, 23156, 12956, 23672, 42008, 37792, 38876, 30488, 27680, 34702, 37724, 37700, 24144, 30744, 33430, 17254, 15982, 23824, 32580, 30826, 27764, 25998, 25276, 34088, 37430, 44478, 20008, 644, 22886, 22138, 29482, 17160, 7916, 10258, 31542, 45500, 30340, 40610, 44368, 40436, 42186, 40796, 42354, 40068, 44188, 31620, 22922, 30236, 29612, 35964, 39748, 44034, 48606, 16968, 0, 1426, 0, 0, 9000, 23318, 24480, 26412, 25508, 26666, 28056, 27802, 27970, 21838, 21334, 26970, 24896, 23558, 24020, 20470, 27552, 38308, 49750, 29282, 30626, 23916, 12312, 24090, 13554, 16664, 15106, 15364, 16258, 13998, 18626, 5488, 7354, 25062, 23756, 27424, 27260, 28504, 29022, 29816, 30312, 30598, 31334, 28464, 33450, 41258, 46798, 37594, 27380, 41212, 35048, 28672, 31848, 24190, 22116, 31060, 24336, 24306, 28570, 20886, 18812, 13700, 16042, 25808, 33848, 30116, 24432, 21536, 26092, 30022, 28756, 29612, 28696, 30038, 27666, 33284, 27034, 24380, 27568, 27250, 27278, 33170, 34224, 19544, 18886, 18650, 17960, 16260, 18472, 19970, 14968, 16106, 15416, 19116, 32604, 29714, 24634, 22340, 22428, 40310, 40172, 48342, 18536, 3034, 10680, 5502, 21160, 24038, 23970, 34548, 45668, 41282, 43618, 41652, 42576, 42038, 42488, 41836, 43056, 40270, 42454, 33116, 34026, 26788, 23936, 37226, 31974, 30730, 34778, 38950, 44466, 32350, 17456, 23154, 26246, 27942, 27854, 29406, 29254, 27554, 27024, 22768, 25872, 21524, 30616, 43934, 36350, 44236, 26794, 26238, 36050, 33654, 36982, 35536, 36548, 37232, 27656, 18322, 21172, 19738, 20540, 20054, 20484, 19064, 16014, 21628, 32212, 23610, 16982, 14274, 25426, 29132, 32980, 41642, 37150, 44260, 24712, 27594, 29916, 21472, 28106, 27244, 19216, 28946, 26858, 12160, 18994, 20246, 18230, 19298, 20050, 14466, 16800, 17318, 19478, 25006, 21488, 19524, 24356, 30006, 34926, 35056, 35310, 34992, 35470, 34666, 36240, 30754, 23446, 26394, 24552, 25472, 17994, 9102, 14616, 18170, 21260, 19838, 19330, 14558, 8824, 2774, 2, 1150, 30670, 48138, 45808, 32380, 19936, 28680, 26836, 26868, 21920, 19890, 23136, 24234, 18320, 16832, 17964, 16606, 18520, 25936, 19628, 14238, 13702, 11074, 11418, 12436, 9672, 15412, 868, 16980, 42068, 39372, 31084, 9466, 30904, 35454, 28680, 27418, 17678, 28324, 36306, 24350, 13748, 23764, 30792, 32846, 28650, 25968, 31526, 34304, 41104, 35546, 45814, 17714, 2004, 17792, 25918, 6160, 19164, 52746, 40736, 40018, 34116, 40230, 38772, 33498, 31310, 31336, 31172, 31432, 30990, 31884, 28450, 23496, 31546, 38718, 37284, 41152, 42668, 45800, 42522, 49754, 22266, 0, 4002, 1182, 12718, 21066, 23036, 23270, 24504, 25590, 22802, 21572, 22538, 18902, 19250, 19824, 20774, 10922, 21314, 43168, 42440, 45272, 48908, 40784, 48390, 22344, 0, 2566, 0, 3022, 1606, 1992, 2386, 1004, 6502, 16666, 21410, 23094, 23534, 24850, 24328, 25976, 26022, 29248, 24482, 31148, 10384, 17678, 47038, 33374, 37890, 30042, 34062, 34530, 22016, 35674, 24508, 13520, 17004, 20564, 22610, 14552, 15534, 14226, 18594, 30330, 35780, 35818, 34536, 35664, 27492, 23436, 27752, 26236, 26656, 27150, 25518, 29086, 19622, 25816, 30110, 32048, 36134, 40448, 20312, 23756, 28102, 8020, 29566, 33350, 30384, 27500, 12522, 9814, 8710, 18274, 36788, 26616, 19666, 26684, 25558, 33814, 42146, 48994, 22642, 0, 4214, 0, 8432, 3164, 21520, 46424, 38716, 43246, 41690, 38090, 34806, 35688, 35428, 35298, 35792, 34724, 37604, 35578, 31286, 35408, 26290, 24538, 34298, 29848, 35824, 38008, 46180, 20368, 5280, 23264, 20094, 24328, 23324, 25588, 24324, 24480, 22054, 23712, 11830, 27886, 46160, 36440, 34700, 33740, 34976, 27620, 19644, 23698, 23412, 18766, 16992, 11110, 17468, 21760, 21684, 21860, 21766, 21778, 21874, 21528, 23544, 30760, 34584, 32020, 32234, 23814, 25582, 38536, 29520, 32952, 36870, 33324, 33326, 34676, 25856, 26184, 22598, 25392, 27404, 7956, 30424, 19660, 8324, 27172, 8222, 8222, 1944, 1757, 595, 5963, 13017, 13757, 16804, 14424, 11554, 13510, 13542, 13740, 13924, 13926, 14091, 14066, 14281, 14029, 14728, 15367, 15261, 15713, 15525, 15017, 15251, 15222, 15455, 15271, 16420, 16927, 17514, 19850, 19030, 17854, 17603, 16132, 15269, 15457, 15447, 15307, 15650, 14909, 17379, 19681, 18393, 17798, 17256, 17304, 17309, 17592, 17477, 17708, 18043, 18286, 18699, 18942, 19676, 20151, 20273, 20595, 20625, 20698, 21276, 21676, 21936, 22269, 22586, 22875, 23005, 23309, 23216, 23362, 23453, 23467, 23513, 23751, 23883, 24304, 25176, 25520, 25586, 25559, 25596, 25532, 25649, 25418, 26111, 26356, 25819, 25759, 25301, 24840, 24857, 24749, 23890, 23146, 22501, 21985, 21552, 21403, 20239, 19231, 18846, 18459, 16458, 14107, 12565, 11035, 6228, 2401, 2569, 2468, 2508, 5380, 9627, 10811, 11401, 11774, 11978, 12332, 12254, 12137, 12152, 12315, 12492, 12438, 12462, 12445, 12465, 12443, 12217, 10260, 10237, 11103, 13978, 16804, 16979, 18393, 18983, 19343, 18502, 18639, 14378, 11402, 12684, 12367, 12968, 13085, 13474, 13598, 13760, 13834, 13892, 13927, 13625, 13523, 13415, 13341, 13145, 12084, 10813, 9350, 6838, 7734, 12272, 16340, 18349, 19838, 20769, 20533, 20585, 20673, 20414, 20989, 18985, 16489, 16464, 15763, 15867, 15762, 15546, 15254, 15008, 14855, 15329, 14492, 17711, 21483, 21613, 22296, 22248, 22091, 21950, 21659, 21052, 20522, 19794, 19201, 17720, 18091, 14272, 10899, 12153, 12083, 12476, 12362, 12175, 12618, 12912, 12784, 13038, 13399, 13646, 13564, 13621, 13559, 13650, 13487, 13967, 14124, 13504, 13382, 12731, 12222, 12066, 11312, 12054, 8619, 6020, 7833, 7531, 7350, 7301, 6294, 10563, 16041, 17405, 19309, 20032, 19568, 19489, 20158, 20772, 20379, 20165, 20271, 19784, 19680, 20353, 21589, 22529, 23136, 23474, 23743, 24058, 23856, 23463, 23687, 23396, 23864, 23048, 24652, 19150, 11967, 13008, 10820, 14370, 18261, 17849, 18713, 18474, 18495, 18439, 18189, 17986, 18202, 18301, 18887, 19415, 19287, 19400, 19473, 19305, 19745, 20111, 20172, 20468, 20473, 21038, 20929, 20147, 19902, 19989, 20324, 20479, 20649, 21125, 21389, 21403, 21431, 21497, 21538, 21398, 21689, 21139, 22244, 18651, 15278, 16383, 16065, 16955, 16475, 13512, 12098, 12776, 13151, 13879, 14031, 14580, 15183, 15246, 13697, 13283, 10186, 8608, 7709, 4340, 4026, 4065, 4283, 4522, 4269, 5380, 8640, 10877, 12240, 13819, 14573, 14502, 14197, 14230, 14272, 14771, 15437, 15416, 15459, 15423, 15465, 15407, 15503, 15237, 15212, 15741, 15004, 15362, 11808, 9274, 11215, 11361, 11948, 12161, 12484, 11968, 13688, 16369, 15914, 17060, 16789, 14498, 13168, 14609, 15942, 15941, 10131, 6067, 7647, 7507, 8582, 9394, 8922, 11063, 14464, 15531, 16799, 17496, 18084, 17950, 18622, 19100, 18962, 19031, 18990, 19015, 18994, 19060, 19233, 19059, 18955, 19226, 19090, 19491, 19684, 20455, 20900, 20785, 21092, 21438, 20454, 20085, 17045, 16518, 19859, 19429, 19507, 18715, 18672, 16909, 14984, 14094, 12310, 13618, 17497, 13713, 10426, 12073, 11908, 12548, 12967, 13639, 13590, 13625, 12958, 12563, 12621, 12677, 12497, 12915, 11446, 9715, 9856, 9960, 9701, 9678, 5274, 1782, 3692, 3494, 6156, 8698, 8932, 8941, 8483, 9434, 9919, 10483, 12319, 13613, 13738, 14981, 16362, 18504, 15976, 13608, 15398, 14594, 16789, 19165, 19240, 19482, 19894, 20401, 20534, 20509, 20415, 19944, 19130, 18934, 18864, 19079, 18645, 19532, 16644, 14062, 15250, 15364, 15727, 16002, 17117, 17154, 17886, 18197, 18424, 19487, 19913, 20497, 20851, 20947, 21223, 21257, 20970, 21459, 21607, 21338, 21140, 21055, 21457, 20294, 19601, 20014, 20207, 20187, 20400, 20191, 19472, 19212, 18746, 18551, 18337, 18394, 18379, 18167, 18258, 18187, 18270, 18135, 18554, 18950, 18626, 18624, 17994, 16816, 16686, 17098, 17276, 17557, 17626, 17794, 18039, 18293, 18498, 18127, 18198, 18432, 17617, 14862, 14528, 14718, 13846, 14351, 14584, 14691, 14503, 14327, 14592, 14636, 10953, 9782, 10147, 13388, 15631, 15048, 17117, 17061, 17819, 18344, 18193, 18265, 18240, 18234, 18019, 15800, 14669, 14862, 14560, 14775, 15001, 14723, 14252, 14357, 14264, 14310, 14153, 14164, 14362, 14294, 14458, 14023, 14511, 12151, 11789, 13578, 11886, 11826, 11855, 11795, 11637, 11548, 11057, 10706, 11783, 11850, 11771, 11740, 13079, 14715, 14069, 16323, 17977, 17445, 17830, 17406, 18028, 16892, 20428, 23288, 21754, 22183, 21334, 19097, 17904, 18217, 16241, 15403, 15757, 15814, 16138, 16027, 16732, 17536, 18204, 19008, 18841, 19123, 19405, 19370, 18841, 18772, 19100, 19036, 19108, 18525, 17281, 15165, 14595, 12770, 14350, 17764, 18038, 19331, 19579, 20371, 20761, 20690, 20665, 20786, 20521, 21088, 18964, 15817, 18188, 20356, 20532, 20843, 20899, 20986, 20737, 20933, 20275, 19638, 19261, 18383, 18596, 18581, 19005, 19098, 19765, 20279, 20138, 18649, 17429, 18431, 18304, 18649, 18579, 18097, 16895, 15713, 15776, 15825, 16396, 16705, 17224, 17346, 17277, 17567, 17613, 17572, 17669, 17477, 17832, 17124, 19468, 21792, 20157, 19945, 19376, 19377, 19767, 20232, 19547, 17761, 17870, 19058, 19408, 19983, 20604, 20855, 21199, 21406, 22021, 22360, 21672, 20904, 20453, 19651, 19827, 19721, 19307, 16522, 14561, 15028, 14811, 15087, 15069, 15123, 15022, 14870, 14866, 14926, 14945, 14878, 15035, 14729, 15298, 14162, 17902, 21753, 19927, 17933, 13375, 13442, 15341, 15672, 16898, 17146, 17226, 17472, 17733, 18019, 17972, 18081, 18032, 17822, 17559, 17561, 17644, 17726, 17995, 17837, 17997, 17640, 17418, 17578, 19418, 21745, 22206, 23050, 23627, 23639, 23620, 23674, 24034, 24284, 24203, 24292, 24152, 24397, 23953, 24836, 21931, 18822, 19271, 19189, 19824, 19364, 19549, 20348, 18867, 19723, 22223, 21532, 21274, 21367, 21301, 21561, 22028, 22432, 22794, 22604, 22062, 21955, 21575, 21167, 20493, 18945, 18555, 18937, 18942, 19633, 19234, 19709, 20433, 19881, 19815, 19932, 18200, 15760, 15532, 15499, 15538, 15492, 15564, 15420, 15937, 17073, 18790, 19778, 19963, 20289, 20144, 20232, 20153, 20096, 19259, 18335, 18172, 17830, 18580, 20032, 20242, 21074, 21762, 22521, 23018, 23466, 24425, 24354, 24678, 24238, 23670, 23472, 23500, 23491, 23433, 22150, 20727, 20127, 19902, 20601, 21192, 21438, 21327, 21368, 21355, 21352, 21385, 21293, 21607, 21653, 21519, 21449, 24483, 18600, 13080, 15073, 14442, 15163, 14757, 15288, 15645, 15590, 15533, 15567, 15701, 15583, 15774, 16070, 16023, 16882, 16196, 18840, 21862, 22403, 22914, 23223, 24471, 24212, 23926, 23849, 24168, 23503, 22946, 22838, 22744, 22705, 22588, 22650, 22581, 22686, 22506, 22857, 21728, 20791, 21372, 20074, 18739, 18766, 19374, 19498, 20168, 21010, 21269, 22025, 22528, 22718, 22455, 22292, 22559, 22388, 22404, 22557, 22592, 22553, 22540, 22603, 22674, 22522, 22812, 22209, 22844, 18433, 14404, 15874, 15525, 15644, 15417, 15864, 16876, 17836, 18179, 18075, 18161, 18047, 18235, 17867, 19050, 20051, 19399, 18940, 20111, 20483, 22117, 24320, 24080, 24362, 24416, 21392, 17707, 16523, 15805, 16991, 18334, 19147, 19355, 19917, 20824, 21152, 21658, 22138, 22556, 22729, 23022, 23330, 23256, 23245, 23289, 23241, 23243, 23278, 23274, 23274, 23307, 23378, 23356, 23362, 23367, 23349, 23386, 23312, 23567, 23775, 23378, 23345, 23535, 23278, 23381, 20581, 18703, 19698, 19850, 20137, 20221, 20196, 20094, 20185, 20198, 20249, 20214, 20289, 20167, 20049, 19321, 19110, 18123, 18526, 19044, 18707, 19399, 19392, 19659, 19968, 20589, 20926, 21275, 21757, 21956, 22029, 22120, 22109, 22074, 22167, 21978, 22362, 21146, 20093, 20089, 20836, 22679, 23108, 23684, 24049, 24146, 24192, 24165, 24320, 24746, 25014, 24827, 24439, 24297, 24330, 24339, 24454, 23765, 24768, 22278, 19989, 20852, 20378, 20684, 20330, 19542, 19501, 15865, 15234, 18227, 18174, 18923, 19660, 20508, 20160, 19867, 19931, 19935, 19868, 20020, 19693, 20857, 22354, 21465, 21582, 21985, 22114, 21976, 23110, 24355, 24316, 25344, 26039, 26380, 26174, 26022, 25200, 24832, 24000, 23553, 22938, 20207, 19862, 20456, 20659, 20951, 20951, 20872, 20894, 20705, 20533, 20928, 21220, 21422, 21168, 21020, 21254, 20808, 20637, 20697, 20656, 20706, 20628, 20763, 20501, 21341, 22166, 22190, 22548, 22398, 22451, 22101, 21907, 22081, 22202, 21859, 22211, 23494, 23689, 23596, 22738, 22496, 21765, 20397, 21597, 22853, 23512, 23371, 22926, 22983, 23090, 23120, 23739, 24564, 24713, 25532, 25851, 25357, 24666, 23973, 24004, 24143, 24265, 24370, 24280, 24421, 24169, 24685, 22809, 19242, 17056, 17790, 19424, 19798, 20187, 20052, 19650, 18716, 18875, 17626, 16723, 17741, 17993, 19114, 21036, 21872, 22510, 22959, 23034, 23266, 23045, 22303, 21424, 21153, 21298, 21671, 22956, 24588, 24327, 23819, 24314, 24340, 24442, 24453, 24438, 24504, 24251, 24076, 24047, 24197, 23875, 24544, 22337, 20234, 21062, 20800, 20933, 20870, 21073, 21211, 21051, 21125, 21230, 21052, 21104, 20908, 20797, 20777, 20796, 20918, 20398, 21008, 21545, 20153, 16991, 16136, 17163, 17486, 18154, 18254, 18280, 18496, 18591, 18604, 18581, 18537, 18557, 18498, 19093, 21137, 22855, 22906, 23000, 22870, 23076, 22689, 23954, 25329, 24809, 25101, 24995, 25558, 23141, 21326, 22119, 22010, 22185, 22128, 22148, 22121, 21793, 20954, 20904, 21243, 21967, 22705, 21134, 20137, 20589, 20576, 21047, 20637, 20712, 20919, 20873, 20813, 20871, 21137, 21067, 21184, 21364, 21276, 21078, 21080, 20826, 20793, 20771, 20819, 20727, 20914, 20278, 19375, 18840, 18286, 18299, 18162, 18653, 18695, 18749, 18846, 18943, 18680, 18355, 18721, 18621, 18779, 18887, 19084, 19232, 19304, 19661, 19490, 19426, 19111, 20635, 22504, 22332, 22767, 22300, 22428, 20283, 18863, 19739, 19328, 19323, 19041, 17883, 17173, 17460, 17309, 17433, 17287, 17508, 17091, 18504, 20275, 19924, 20902, 21946, 22209, 22187, 22254, 22567, 22947, 23057, 23155, 23508, 23608, 23631, 23517, 23053, 23330, 21934, 20924, 19220, 18694, 20182, 20750, 19455, 18207, 18907, 18640, 18754, 18748, 19061, 18890, 18883, 18783, 19532, 21053, 21007, 20005, 19591, 19708, 19617, 19733, 19546, 19901, 18780, 17794, 18105, 18008, 18467, 18132, 17971, 18086, 17995, 18207, 18041, 17709, 17333, 16761, 16168, 17069, 17927, 17542, 18422, 19384, 19539, 19991, 20322, 21070, 21710, 21666, 21880, 22214, 22582, 22797, 22669, 22435, 22064, 21702, 21716, 21713, 21707, 21894, 22033, 22025, 21966, 22114, 21820, 22407, 20637, 19666, 19676, 18802, 20597, 21305, 21482, 21531, 21557, 21457, 21359, 21499, 21393, 21350, 19920, 18926, 18706, 18423, 18417, 18086, 18360, 18627, 18477, 18963, 15988, 14044, 15261, 14893, 15525, 15560, 16261, 16868, 16708, 17522, 18387, 18918, 19415, 19597, 19500, 19537, 19521, 19523, 19534, 19503, 19623, 19817, 19682, 19356, 18747, 18631, 18987, 18979, 19070, 19221, 19241, 19229, 19256, 19451, 19466, 19495, 19585, 19483, 19491, 19090, 19051, 18624, 19923, 21273, 20986, 19798, 18072, 16715, 15949, 15592, 15945, 13186, 10746, 11554, 11263, 11585, 11592, 11473, 11313, 11319, 11402, 11204, 11592, 10817, 13218, 15184, 15600, 15984, 12279, 14424, 16456, 16896, 15142, 14984, 18173, 18721, 20667, 21928, 22661, 23012, 23339, 23189, 23412, 22630, 21029, 18837, 17716, 18310, 18238, 18228, 18136, 18340, 18817, 19041, 19013, 19159, 19515, 19117, 19610, 16762, 13032, 16380, 18372, 17866, 18123, 17963, 18075, 17980, 18134, 18015, 17501, 17535, 14746, 13571, 15655, 16217, 16236, 16393, 16848, 16944, 17645, 18562, 18901, 19146, 19317, 19398, 19540, 19590, 19848, 19661, 18775, 18503, 18553, 18565, 18525, 18544, 18492, 18425, 18394, 18398, 18451, 18489, 18083, 18903, 20132, 20470, 20737, 20732, 20570, 20955, 20203, 21726, 16744, 11926, 13485, 12780, 13066, 12461, 12647, 12765, 12898, 12881, 13031, 12835, 13169, 12329, 14786, 17330, 17031, 18422, 18626, 18450, 18630, 18293, 18279, 14298, 11964, 14142, 14427, 16391, 18218, 16436, 15107, 16042, 16757, 16738, 17139, 15379, 16501, 19791, 19602, 19867, 19654, 19880, 19559, 20145, 18229, 16127, 16963, 16108, 16995, 13942, 10687, 12016, 10792, 13658, 16442, 16049, 16130, 15764, 15216, 15288, 12452, 9866, 10985, 10218, 12413, 14785, 14680, 14852, 15142, 15604, 16353, 16219, 17127, 18474, 17915, 17748, 17798, 18020, 18358, 18513, 18461, 18693, 18867, 18792, 18877, 18748, 18967, 18544, 19902, 20609, 17617, 16792, 17672, 17735, 17755, 18050, 18145, 18040, 18088, 18071, 17881, 17587, 17167, 17396, 16530, 17260, 13217, 9839, 11460, 11583, 12185, 11954, 12098, 12143, 12241, 12205, 12199, 12147, 12107, 12123, 12401, 12359, 12233, 12330, 12624, 12752, 12685, 12678, 12745, 12593, 12888, 12289, 14297, 16649, 16557, 17060, 17107, 17265, 16761, 16243, 17499, 16616, 15594, 16682, 16878, 17113, 17238, 17302, 17042, 16690, 16840, 16149, 15571, 12149, 9276, 10078, 9680, 10004, 10362, 10432, 10495, 10612, 10663, 10681, 10896, 10569, 11116, 12659, 13363, 13618, 13725, 13649, 13771, 13565, 13925, 13217, 15670, 18934, 17917, 19317, 15551, 11692, 13586, 16701, 18234, 17572, 18034, 18064, 18302, 18196, 18319, 18112, 18105, 17345, 17722, 19419, 20275, 19478, 17371, 16524, 17103, 13644, 11225, 11622, 11357, 9747, 10912, 2440, 4921, 14276, 12209, 14055, 13717, 14251, 13773, 13978, 13846, 13989, 13759, 14208, 12789, 11750, 12072, 12163, 11448, 13346, 8445, 3178, 4653, 3724, 4914, 5078, 5456, 6440, 5541, 8487, 12543, 13314, 14399, 15100, 15612, 16124, 17003, 17421, 17747, 17483, 14454, 12771, 13279, 12934, 13090, 12888, 13196, 13327, 13000, 13118, 12991, 12836, 12815, 12781, 12864, 12703, 13002, 12407, 14315, 15955, 15244, 15633, 15472, 15773, 15694, 15632, 15569, 15992, 16185, 16605, 17280, 17012, 16287, 16861, 13930, 11350, 12129, 12016, 12837, 13269, 13904, 13983, 15018, 16612, 17344, 17780, 17787, 17928, 17938, 17962, 17674, 17257, 17053, 16962, 17011, 16939, 16942, 16904, 16982, 16834, 17136, 16142, 15146, 15285, 15456, 14384, 13539, 13288, 12923, 13571, 14569, 14969, 15259, 15770, 15580, 16002, 16428, 16112, 16658, 14104, 11759, 12361, 12210, 11834, 11473, 11749, 11972, 13607, 14369, 14924, 15198, 14649, 14518, 14376, 15709, 17184, 17594, 17609, 17446, 17543, 17679, 17486, 17849, 17171, 18516, 14313, 10806, 10291, 10125, 12996, 11635, 11593, 12341, 12370, 12080, 11344, 9099, 5921, 2340, 8128, 13404, 12579, 13628, 13649, 13544, 13179, 13010, 12733, 12375, 12384, 11307, 10385, 10978, 11891, 12671, 13713, 14424, 14516, 15401, 15238, 15776, 16130, 16306, 17223, 17387, 17407, 17342, 17467, 17212, 18087, 19073, 18604, 18675, 18302, 17361, 17473, 17072, 18212, 14061, 12680, 11272, 8334, 11162, 11339, 12014, 12240, 12351, 12323, 11068, 9186, 5925, 5632, 9754, 11712, 11812, 12530, 11737, 15201, 15201, 124, 0, 0, 105, 297, 88, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 123, 0, 435, 0, 3511, 7932, 6807, 7197, 7209, 4044, 78, 111, 0, 33, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 2, 458, 4456, 6739, 6191, 6327, 6487, 5969, 7140, 3171, 0, 393, 0, 112, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 62, 0, 658, 2445, 3294, 3721, 3948, 4379, 4354, 5080, 5773, 5555, 5675, 5596, 5658, 5581, 5935, 6868, 5327, 3995, 1539, 0, 185, 0, 45, 0, 0, 23, 0, 398, 1859, 2656, 3378, 4583, 5408, 4764, 4512, 4506, 3969, 4072, 3738, 2949, 1813, 1606, 2087, 745, 0, 80, 0, 23, 0, 5, 0, 0, 0, 0, 0, 0, 2, 0, 12, 0, 47, 0, 403, 1165, 2070, 3418, 4149, 4522, 4577, 4582, 4490, 4430, 4416, 4476, 4475, 4658, 3768, 4201, 7696, 8544, 7995, 8528, 8681, 8694, 8391, 8270, 8155, 10150, 7954, 4265, 4625, 4401, 3870, 2259, 874, 627, 721, 698, 697, 723, 661, 793, 352, 0, 43, 0, 8, 0, 174, 1543, 2232, 2822, 3307, 3008, 1118, 0, 130, 0, 37, 0, 19, 0, 49, 0, 400, 1194, 2956, 5992, 7204, 8173, 8515, 11266, 11321, 9398, 10461, 11217, 10793, 8250, 6697, 5900, 5740, 5756, 5777, 5714, 5842, 5575, 6558, 8318, 9074, 10066, 10174, 10386, 10808, 10665, 10872, 10254, 9346, 8500, 8031, 8395, 8343, 7873, 7708, 5966, 6145, 2710, 0, 339, 0, 96, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 82, 0, 284, 0, 2606, 7645, 8240, 9280, 9949, 10463, 10874, 10900, 10936, 11061, 10885, 10648, 10388, 10161, 9980, 9628, 9054, 7967, 6486, 3325, 1134, 376, 0, 152, 2416, 4806, 4948, 5414, 6150, 6849, 7113, 7252, 7511, 7748, 7255, 6908, 7082, 6851, 7236, 6551, 7892, 3514, 0, 533, 0, 471, 0, 2844, 6488, 5651, 7023, 7711, 9000, 9283, 9405, 8374, 7851, 7333, 8268, 3583, 0, 441, 0, 150, 0, 150, 0, 433, 0, 3685, 9386, 8588, 9277, 9432, 10047, 9608, 10422, 11641, 11219, 11090, 11186, 10977, 11384, 10635, 12121, 7221, 2068, 4175, 4218, 6419, 2635, 0, 316, 0, 95, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 37, 0, 125, 0, 2570, 7235, 8978, 9456, 9167, 8963, 9121, 8854, 9335, 8459, 10195, 4509, 0, 560, 0, 160, 0, 32, 0, 0, 1, 0, 1, 0, 0, 0, 222, 1718, 1283, 524, 770, 2173, 3180, 4297, 4746, 4913, 6560, 7137, 6580, 5356, 5665, 5379, 5099, 5258, 5406, 5322, 5225, 5384, 5219, 5053, 5158, 5000, 5276, 4779, 5762, 2548, 0, 316, 0, 90, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 20, 0, 65, 0, 640, 1814, 620, 0, 62, 0, 15, 0, 0, 10, 0, 41, 0, 869, 5027, 7568, 7862, 8228, 8036, 8231, 7955, 8415, 7529, 10401, 13235, 12370, 13784, 13240, 12693, 11994, 11700, 11984, 12904, 14919, 14855, 14740, 15222, 14501, 13947, 13759, 13718, 12258, 11430, 4143, 0, 2206, 3105, 3664, 5481, 7586, 9536, 11596, 12356, 13833, 14281, 14880, 15651, 15956, 15594, 16771, 14345, 11749, 12679, 11956, 12813, 11502, 13935, 6414, 1401, 7305, 7387, 7734, 5921, 3179, 1439, 1531, 3267, 4194, 4333, 4881, 6017, 5644, 3271, 2032, 2133, 1059, 1110, 2786, 3486, 3891, 3892, 4487, 6066, 7675, 7826, 8077, 8735, 9596, 9523, 10528, 11370, 11457, 11664, 11653, 11305, 10981, 11051, 11067, 10967, 11186, 10725, 12290, 14089, 13802, 14532, 15030, 15550, 15799, 16076, 16168, 15456, 14870, 14593, 14463, 14091, 12571, 9258, 8961, 3602, 0, 430, 0, 111, 0, 0, 77, 0, 589, 580, 0, 44, 33, 0, 277, 0, 2552, 7163, 8006, 8878, 8713, 8780, 8826, 8644, 9031, 8204, 8918, 3716, 0, 451, 0, 128, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 64, 807, 2109, 3209, 4494, 6173, 7218, 7514, 7703, 8117, 8785, 9174, 8274, 7767, 8016, 8026, 7754, 7545, 8063, 7962, 8110, 7466, 6897, 6914, 7172, 6550, 7880, 3457, 0, 322, 0, 0, 1837, 5464, 6237, 5849, 7262, 3296, 0, 412, 0, 117, 0, 23, 0, 0, 0, 0, 0, 0, 13, 0, 61, 0, 208, 0, 2141, 7274, 7890, 7634, 8222, 8555, 8847, 8727, 9048, 9649, 9636, 9682, 9625, 9711, 9600, 9112, 3039, 0, 367, 0, 575, 2892, 8783, 10493, 8101, 7025, 6084, 5905, 7372, 9685, 13956, 12301, 9076, 10352, 10033, 10337, 9853, 9947, 8992, 8966, 3406, 0, 396, 0, 113, 0, 15, 4, 0, 85, 0, 292, 0, 3859, 7549, 6538, 6895, 6963, 6387, 8709, 11077, 10267, 10585, 10324, 9929, 8914, 8064, 7213, 7028, 8120, 9046, 9477, 9641, 10319, 11393, 11787, 11738, 11979, 11752, 11269, 11462, 10928, 9628, 7799, 2337, 0, 236, 0, 68, 0, 14, 0, 0, 0, 0, 0, 0, 28, 0, 141, 0, 496, 0, 3955, 8800, 7564, 9164, 8591, 7943, 7071, 6519, 6442, 5254, 4210, 3797, 3896, 3984, 4443, 5251, 5140, 5408, 5665, 5959, 6162, 5022, 4442, 5124, 6083, 6833, 6746, 7411, 7373, 7029, 7274, 7521, 7826, 7518, 7434, 6655, 5808, 5859, 5757, 5869, 5693, 6002, 5441, 6557, 2901, 0, 360, 0, 101, 0, 20, 0, 10, 0, 29, 122, 2109, 4024, 4350, 3911, 2495, 671, 0, 65, 0, 51, 33, 826, 0, 4585, 8254, 8759, 3756, 0, 0, 2476, 6775, 6175, 7097, 6127, 6080, 6551, 6565, 6660, 6478, 6796, 6223, 7363, 3456, 0, 1723, 3367, 6482, 7965, 9608, 10751, 8925, 6838, 5117, 5210, 5147, 5003, 5563, 5204, 6824, 10001, 6843, 3923, 3972, 3708, 3939, 3756, 3489, 3359, 2742, 2889, 3212, 3942, 6644, 9361, 10599, 11905, 13418, 13760, 14259, 14571, 14463, 14531, 14461, 14560, 14406, 14685, 13766, 12486, 12468, 10858, 11545, 4543, 0, 536, 0, 154, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 67, 0, 234, 0, 1905, 4336, 3618, 4174, 4754, 5444, 5691, 5909, 5867, 6046, 6549, 6999, 6974, 7196, 7461, 7523, 7745, 8010, 8456, 8799, 9188, 9248, 9309, 9464, 10039, 9672, 9912, 9046, 8961, 4079, 0, 2060, 3228, 4282, 5023, 6094, 6547, 2844, 333, 1005, 745, 751, 1001, 357, 2302, 2620, 2297, 2647, 1288, 1625, 1503, 3193, 6373, 9824, 11799, 12555, 12862, 13183, 13104, 12858, 8465, 5642, 6626, 6481, 6904, 6836, 6851, 6841, 6893, 6831, 6869, 6803, 6515, 2868, 1950, 3974, 5591, 6970, 6686, 7392, 7693, 7898, 7881, 7907, 7862, 7944, 7780, 8145, 6607, 2193, 0, 3358, 8507, 9474, 9521, 10813, 4701, 0, 494, 0, 53, 91, 0, 577, 0, 5057, 13228, 13495, 15785, 16168, 16647, 16709, 16471, 16696, 16410, 16230, 13722, 12040, 12831, 12892, 13362, 13219, 13234, 13468, 13749, 13973, 14000, 13999, 14000, 13998, 14002, 14001, 14016, 13976, 13470, 12892, 12307, 11555, 9808, 2914, 0, 287, 0, 83, 0, 32, 0, 28, 401, 5043, 8932, 8651, 9872, 12978, 14752, 15132, 13182, 9919, 11468, 4590, 0, 467, 0, 0, 1478, 8865, 13596, 14456, 15249, 14989, 14865, 14958, 14777, 15114, 14493, 15721, 11702, 7706, 9023, 8415, 8741, 8628, 8693, 8820, 9267, 9248, 9166, 9249, 9503, 9497, 9792, 9630, 9598, 7169, 5075, 5113, 4431, 4826, 4658, 4939, 5452, 7431, 9226, 8445, 7936, 6392, 1673, 0, 149, 0, 43, 0, 9, 0, 14, 0, 73, 0, 257, 0, 2091, 4875, 4315, 4938, 4623, 5226, 6102, 6861, 7413, 7638, 7892, 8299, 7696, 8009, 6504, 9529, 13161, 10348, 10103, 10471, 10509, 10790, 10902, 11229, 11180, 11818, 13114, 14093, 14758, 14826, 14266, 13771, 13808, 13665, 13582, 13413, 13764, 12974, 12269, 12461, 12397, 12375, 12494, 12216, 13251, 15047, 15146, 15699, 14948, 17177, 10903, 5952, 3409, 0, 483, 0, 75, 24, 0, 1667, 3875, 3915, 4076, 4203, 4337, 4019, 4491, 2350, 0, 684, 0, 4433, 10747, 9716, 10614, 10109, 10113, 10205, 10218, 10072, 10157, 10295, 10251, 10266, 10273, 10242, 10309, 10171, 10585, 10722, 10225, 9390, 8599, 8565, 8902, 8459, 10676, 6931, 2813, 3797, 2475, 5205, 3245, 4195, 6894, 4578, 4463, 5022, 5921, 5431, 5690, 6055, 5979, 5720, 5049, 5544, 5768, 4484, 3808, 4246, 4888, 5784, 5942, 6095, 5051, 1437, 0, 315, 150, 238, 195, 205, 249, 357, 575, 648, 723, 699, 600, 760, 724, 232, 0, 22, 0, 5, 0, 0, 42, 0, 199, 0, 923, 0, 6006, 12989, 12973, 14862, 13925, 15503, 17106, 17518, 17501, 16841, 17250, 16906, 14867, 13620, 13672, 13170, 13085, 12798, 13440, 12207, 14697, 6506, 0, 808, 0, 230, 0, 37, 0, 0, 48, 224, 3550, 5777, 5431, 5776, 6098, 6868, 7370, 6975, 7978, 4302, 0, 210, 0, 64, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 167, 0, 597, 0, 4484, 8593, 6060, 3677, 0, 222, 0, 285, 2330, 3978, 3876, 4734, 5598, 6114, 6489, 6373, 6634, 5489, 4333, 1605, 0, 189, 0, 52, 0, 9, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 17, 0, 166, 247, 394, 38, 733, 0, 3974, 8823, 7479, 8386, 6309, 4972, 2269, 0, 124, 0, 35, 0, 4, 0, 0, 13, 0, 66, 0, 228, 0, 2000, 5327, 5080, 6265, 7180, 7495, 7964, 8242, 8294, 8527, 8512, 8691, 8578, 7895, 2896, 0, 234, 702, 1510, 1232, 1362, 1312, 1308, 1412, 1508, 1413, 1245, 1049, 786, 196, 0, 17, 0, 4, 0, 1, 0, 0, 16, 0, 81, 0, 285, 0, 2496, 6679, 6707, 7541, 8805, 9578, 10981, 10290, 13986, 14145, 10490, 11790, 11370, 11759, 11961, 11888, 11450, 11506, 11468, 11489, 11480, 11480, 11483, 11526, 11899, 11957, 11444, 11760, 11369, 12018, 10813, 14807, 19084, 18315, 18360, 18699, 14882, 11855, 13237, 12512, 13163, 13065, 12564, 11740, 11052, 10980, 10817, 10666, 11083, 11187, 10717, 9385, 7705, 5872, 6892, 2965, 0, 361, 0, 103, 0, 21, 0, 0, 9, 0, 48, 0, 173, 0, 1678, 5641, 7772, 8798, 8842, 9364, 9855, 9915, 9898, 9968, 9729, 9432, 9279, 8933, 8289, 8470, 7590, 6317, 5687, 5316, 5582, 5658, 6197, 6507, 7367, 8170, 8764, 9249, 9276, 9531, 9395, 9430, 9449, 9601, 9363, 9090, 9177, 9133, 9163, 9134, 9180, 9055, 8949, 8208, 6341, 1846, 0, 184, 0, 52, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 90, 0, 319, 0, 2746, 7438, 8603, 10299, 10522, 11055, 10812, 11243, 12002, 11657, 11427, 11532, 11383, 11665, 11131, 12121, 10195, 15717, 16133, 11355, 13056, 11459, 11905, 11521, 11241, 11152, 11064, 10901, 10299, 9131, 8570, 8402, 8803, 8571, 8450, 6996, 6006, 5284, 8896, 13476, 13764, 14214, 12544, 3969, 0, 463, 0, 303, 0, 1550, 3771, 4203, 4798, 4425, 4540, 4426, 4524, 4386, 4623, 4186, 5057, 2212, 0, 211, 0, 0, 1134, 4113, 4505, 6145, 7434, 7637, 8408, 8259, 8371, 8653, 8656, 8889, 8858, 8942, 9291, 9308, 9617, 9645, 9806, 10107, 10225, 10020, 9474, 8926, 8345, 7710, 7553, 5345, 4296, 1855, 0, 235, 0, 67, 0, 24, 0, 52, 0, 414, 974, 1855, 2125, 2981, 1503, 0, 125, 193, 486, 604, 1069, 1225, 1238, 1129, 1319, 1247, 1199, 849, 905, 743, 2186, 6059, 6633, 7180, 7200, 6879, 7231, 7226, 7047, 8047, 3462, 0, 421, 0, 112, 0, 161, 193, 97, 313, 0, 662, 0, 4186, 9707, 8675, 9621, 9189, 9545, 9912, 9874, 10493, 9713, 10833, 4503, 0, 545, 0, 156, 0, 31, 0, 0, 0, 0, 0, 16, 0, 78, 0, 272, 0, 2328, 6031, 5733, 6513, 6633, 7600, 7832, 7805, 8090, 7867, 7917, 7983, 7775, 8203, 7336, 9989, 11406, 10002, 10097, 8925, 9389, 9613, 11063, 12275, 12215, 12324, 12512, 13001, 13361, 13799, 13688, 13731, 14114, 14108, 13507, 12479, 11879, 3957, 0, 425, 0, 124, 0, 33, 0, 54, 150, 273, 101, 114, 472, 246, 87, 136, 114, 124, 123, 115, 137, 60, 0, 7, 0, 2, 0, 0, 5, 0, 30, 0, 111, 0, 1039, 3233, 4118, 2790, 2074, 1077, 0, 148, 0, 40, 0, 6, 0, 0, 0, 9, 0, 48, 0, 168, 0, 1441, 3763, 3862, 4389, 4320, 4424, 4283, 4508, 4114, 4885, 2273, 0, 585, 0, 2747, 6719, 6497, 7101, 7524, 8151, 9140, 10173, 10246, 10626, 10695, 10925, 11076, 11123, 11353, 8025, 3473, 2417, 2186, 1837, 2191, 2274, 2074, 1548, 724, 521, 518, 724, 1041, 1081, 1046, 1133, 1248, 1446, 1617, 1569, 1586, 1590, 1564, 1626, 1402, 1109, 1063, 464, 13, 9, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 24, 0, 113, 0, 994, 2744, 4399, 4399, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 124, 0, 437, 0, 4239, 12248, 9920, 9252, 20241, 22046, 17863, 18699, 18449, 17980, 15563, 16451, 18327, 22839, 20936, 17840, 18910, 18506, 18686, 18710, 18462, 19023, 17879, 21260, 22394, 21682, 24015, 23548, 23253, 22360, 18152, 11848, 2966, 13262, 14348, 5486, 8075, 5460, 7671, 6704, 5912, 5018, 5009, 1971, 0, 233, 0, 65, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 606, 7809, 22469, 28150, 26333, 21809, 18597, 18105, 17451, 17987, 19005, 20152, 20954, 21564, 20759, 21522, 21883, 22163, 22471, 22097, 22216, 22037, 23129, 22831, 24079, 25260, 23865, 23948, 23373, 17378, 11932, 17186, 21674, 22358, 15498, 7303, 6537, 5484, 4955, 5144, 4936, 5243, 4729, 5719, 2527, 0, 314, 0, 89, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 58, 0, 208, 0, 2356, 8084, 5539, 0, 5968, 22382, 28137, 28008, 27327, 27556, 23318, 20123, 21743, 20647, 20646, 20279, 20616, 20924, 20590, 20642, 20573, 20661, 20517, 20776, 20269, 21857, 23613, 26082, 30175, 31356, 32357, 31387, 28985, 28455, 22362, 24631, 19596, 12472, 9781, 1650, 845, 0, 134, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 104, 0, 518, 0, 1823, 0, 14479, 31874, 26114, 25040, 19810, 21888, 22298, 21905, 21456, 20983, 20651, 20442, 20539, 21597, 22080, 22324, 22087, 21569, 22682, 22531, 24485, 25485, 22610, 15382, 2937, 63, 2293, 2760, 3142, 3143, 2632, 1678, 2565, 3414, 5292, 3354, 1463, 4076, 4564, 4598, 4479, 4705, 4279, 5144, 2280, 0, 282, 0, 80, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 77, 0, 181, 0, 2864, 10981, 1383, 9033, 28015, 29627, 30961, 30011, 29553, 28923, 29512, 29286, 30142, 31235, 30411, 33383, 27780, 38167, 10923, 13913, 34804, 36781, 12092, 14937, 24006, 0, 5941, 1251, 2639, 3912, 0, 16259, 32427, 23696, 26722, 24566, 22998, 15008, 3130, 490, 335, 0, 55, 0, 15, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 185, 0, 638, 0, 5161, 11464, 8223, 13195, 17736, 24552, 28661, 27285, 28302, 27163, 28975, 23504, 18168, 19495, 18875, 19780, 20512, 21300, 21297, 20612, 21635, 20308, 31945, 16655, 0, 3090, 371, 1862, 2613, 2479, 5234, 0, 14961, 32078, 22912, 23022, 21321, 20049, 19384, 8226, 0, 831, 0, 0, 1990, 5946, 6526, 7343, 7402, 7788, 8023, 7778, 8206, 7431, 8961, 3963, 0, 494, 0, 148, 0, 75, 34, 0, 7, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 59, 0, 288, 0, 1014, 0, 7766, 14688, 8746, 10757, 15106, 19480, 24355, 30231, 30504, 28965, 26209, 21278, 18384, 19162, 18803, 18273, 18747, 19336, 20879, 25816, 29174, 29883, 32595, 29692, 36775, 16223, 0, 5513, 2631, 4524, 3802, 4240, 3815, 4504, 3210, 5658, 885, 14339, 13100, 0, 3628, 943, 2095, 1164, 1305, 960, 1095, 446, 0, 53, 0, 15, 0, 2, 0, 3, 0, 28, 0, 56, 64, 1874, 2642, 686, 6873, 4398, 0, 603, 0, 176, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 129, 0, 475, 0, 4263, 12150, 12992, 6282, 6731, 20661, 26174, 26028, 20846, 17644, 18733, 18497, 18503, 18202, 18296, 18274, 18242, 18337, 18138, 18766, 19260, 19328, 19609, 19334, 19321, 19123, 19211, 20308, 23524, 25193, 23218, 27141, 31474, 30832, 25766, 23295, 13955, 2113, 9733, 13728, 11139, 10376, 6020, 3218, 4662, 5668, 5755, 5722, 6029, 5631, 6181, 2614, 0, 319, 0, 91, 0, 34, 0, 82, 0, 291, 0, 1912, 1912, 0, 291, 0, 82, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 219, 0, 746, 0, 6215, 15153, 11736, 13988, 13393, 19182, 21657, 17989, 19451, 18656, 19504, 19699, 19457, 19717, 19983, 20034, 19927, 20314, 20406, 19623, 19117, 18853, 19132, 20596, 23375, 24067, 23216, 24190, 23175, 20544, 8113, 3906, 6828, 8857, 8444, 4507, 5896, 5189, 5578, 5356, 5528, 5139, 4406, 4496, 3931, 4822, 2152, 0, 268, 0, 76, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 153, 0, 515, 0, 4447, 9781, 2472, 6553, 19948, 20340, 17227, 18368, 17419, 17612, 17058, 15978, 16208, 16736, 17425, 17836, 17732, 17746, 17817, 17632, 17987, 17457, 21193, 23856, 22558, 23395, 23504, 23500, 24146, 23090, 21187, 21262, 21729, 20999, 19450, 18084, 16974, 9686, 1142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 237, 0, 843, 0, 5523, 5523, 0, 843, 0, 237, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 26, 0, 99, 0, 896, 2699, 3846, 4683, 4932, 3028, 1476, 1612, 1144, 459, 0, 55, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 143, 0, 595, 506, 10991, 6940, 5871, 22813, 26358, 28979, 30221, 30569, 30019, 30917, 29796, 31757, 27775, 34367, 16216, 0, 3261, 148, 2453, 1635, 2230, 2134, 2616, 2913, 2808, 2899, 2724, 3107, 2280, 4277, 2489, 5371, 0, 17106, 33399, 21932, 22252, 19453, 20460, 18558, 18061, 8598, 0, 11298, 11606, 466, 5441, 3834, 4658, 4547, 2198, 0, 263, 0, 94, 0, 139, 0, 442, 0, 6334, 9465, 7531, 3764, 0, 514, 0, 137, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 117, 116, 4348, 8412, 14601, 17988, 11885, 14834, 18350, 17324, 17815, 17597, 17588, 18001, 18326, 19078, 19648, 20274, 21905, 23358, 25047, 26046, 20808, 31913, 15811, 0, 3861, 1523, 3453, 3511, 4747, 4288, 3865, 5097, 3600, 5466, 0, 16014, 34913, 25896, 27928, 24602, 24303, 21970, 16328, 4717, 0, 635, 0, 277, 111, 210, 218, 213, 228, 219, 222, 173, 0, 236, 0, 1593, 2505, 1090, 668, 0, 103, 0, 24, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 94, 0, 264, 401, 10579, 12674, 453, 4523, 18150, 19500, 16957, 18742, 18207, 18635, 19083, 18971, 19029, 19254, 19416, 19150, 19723, 20756, 20509, 20070, 20184, 20885, 20397, 20055, 20746, 20887, 23188, 23010, 21463, 22164, 21485, 22421, 20887, 23836, 14036, 3215, 7046, 2119, 436, 1652, 1282, 1697, 515, 0, 53, 0, 18, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 88, 0, 325, 576, 10956, 5357, 6690, 25554, 28969, 29030, 26646, 21996, 18949, 19715, 19510, 19329, 19955, 18506, 23458, 29055, 28660, 24857, 20017, 21017, 20231, 19475, 19522, 20243, 20396, 22393, 24952, 22524, 26563, 31820, 30647, 22125, 24273, 16573, 5324, 7400, 2352, 1784, 1765, 789, 0, 77, 0, 22, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 53, 0, 273, 0, 984, 0, 7642, 15647, 13309, 5261, 0, 0, 7563, 19118, 16810, 18511, 17772, 17617, 17559, 18518, 19444, 20033, 19683, 19533, 19383, 19273, 19306, 18940, 20033, 20707, 21379, 20789, 22264, 22425, 22118, 12791, 20348, 32757, 28481, 27806, 25247, 26485, 25353, 26895, 24319, 29332, 12970, 0, 1611, 0, 461, 0, 93, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 11, 0, 0, 0, 1826, 11473, 6887, 3672, 21560, 28364, 26502, 21768, 17984, 18525, 18569, 18529, 19187, 20306, 19845, 19819, 19780, 19832, 19747, 19895, 19616, 20375, 19968, 18378, 18838, 19554, 22903, 25192, 23039, 20555, 26045, 21412, 20911, 23777, 22679, 14452, 4626, 6475, 4235, 4108, 3722, 2382, 198, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 194, 0, 651, 0, 6360, 19832, 18172, 16434, 17343, 17449, 18352, 18566, 18144, 18477, 19066, 19220, 19857, 20511, 20645, 20639, 20165, 19951, 19275, 18922, 18992, 19531, 19551, 21877, 22257, 26200, 11610, 0, 4733, 4355, 3267, 3697, 3597, 2713, 1926, 1828, 1425, 1588, 1528, 1527, 1587, 1448, 1741, 771, 0, 95, 0, 27, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 100, 0, 418, 0, 3908, 10710, 10259, 0, 12165, 27727, 23590, 21186, 16674, 19206, 18378, 19183, 18847, 20230, 21406, 21117, 21304, 20782, 20713, 20568, 20670, 20509, 20068, 20187, 20190, 20077, 20373, 19695, 22150, 26648, 31380, 28003, 23212, 10129, 2504, 6659, 5646, 4314, 11028, 24346, 16333, 7993, 7903, 2952, 165, 12, 0, 14, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2882, 2587, 2333, 865, 2768, 0, 11249, 24698, 23969, 27646, 27262, 27823, 27794, 28141, 28077, 28059, 28528, 27733, 27692, 27083, 27310, 25572, 23862, 9335, 0, 822, 0, 237, 0, 46, 0, 0, 0, 0, 1, 0, 5, 0, 18, 0, 193, 699, 965, 1930, 2485, 2596, 2777, 2809, 2645, 2590, 2891, 2897, 2970, 3129, 3159, 3195, 3141, 2970, 2763, 2923, 2259, 1318, 1386, 1213, 1192, 845, 161, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 6, 0, 72, 349, 955, 1382, 1458, 1734, 1928, 2319, 2361, 2328, 2869, 3053, 3189, 3315, 3274, 3297, 3280, 3297, 3278, 3250, 2716, 2508, 2713, 2274, 2234, 2136, 1931, 1755, 1522, 1648, 1596, 1670, 1767, 1890, 2364, 2926, 3290, 3424, 3357, 3271, 3380, 3414, 3162, 3385, 3638, 3480, 3359, 3132, 3144, 3114, 2978, 2362, 2299, 1067, 0, 94, 0, 27, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 15, 0, 157, 518, 698, 859, 1082, 1135, 1376, 2000, 2305, 2565, 2840, 2934, 2986, 2993, 3277, 2887, 3894, 4376, 4690, 5008, 5362, 6854, 6985, 6856, 7206, 6495, 7828, 5145, 14270, 25679, 24594, 26534, 25919, 26066, 26546, 23517, 26378, 11588, 0, 2121, 281, 1290, 873, 1305, 1215, 1606, 1871, 2135, 2192, 2318, 2437, 3555, 4470, 4259, 4641, 4788, 5033, 5088, 5210, 5183, 4972, 5146, 5109, 4968, 4593, 4240, 4305, 4172, 4403, 3988, 4808, 2127, 0, 264, 0, 75, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 171, 0, 626, 0, 8940, 19916, 23558, 26187, 24937, 26640, 26242, 26980, 27511, 27510, 27453, 27589, 27398, 27157, 25850, 22939, 20159, 8187, 1092, 2459, 1697, 2000, 1873, 1920, 2827, 4121, 4630, 5204, 5222, 5113, 4960, 4950, 4987, 5131, 5208, 5109, 5087, 5098, 5078, 5116, 5041, 5294, 5603, 5562, 5744, 5431, 5139, 5103, 4989, 4905, 4766, 4552, 3999, 1266, 0, 132, 0, 38, 0, 5, 0, 22, 0, 124, 0, 419, 0, 6794, 14822, 14170, 15917, 14787, 17283, 7194, 0, 878, 0, 251, 0, 56, 0, 28, 0, 102, 0, 841, 2033, 2201, 2623, 2814, 1561, 29, 43, 0, 13, 0, 0, 0, 0, 10, 0, 36, 0, 440, 1858, 2758, 3108, 3389, 3683, 3829, 4074, 4316, 4518, 4607, 4515, 4552, 4461, 4412, 4580, 4712, 4789, 4949, 4920, 4817, 4852, 4833, 4845, 4836, 4846, 4824, 4731, 4176, 3094, 2343, 1739, 1547, 1676, 2258, 3007, 3279, 3477, 3550, 3792, 4279, 4539, 4875, 5031, 4758, 4643, 4474, 4268, 4343, 4386, 4284, 4105, 3813, 1286, 0, 139, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 0, 29, 0, 266, 710, 419, 588, 1028, 1315, 1084, 978, 436, 0, 55, 0, 15, 0, 2, 0, 11, 0, 44, 0, 145, 0, 2269, 11006, 14808, 16077, 18963, 18410, 18817, 14192, 4343, 842, 995, 927, 963, 977, 893, 1085, 684, 2026, 3417, 3203, 3684, 3989, 4431, 4580, 4828, 4925, 4851, 4793, 5108, 5259, 5336, 5706, 5902, 6018, 5985, 5662, 5428, 5194, 5120, 4867, 4640, 4778, 4475, 4272, 4253, 3891, 4047, 1530, 0, 176, 0, 51, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 170, 0, 476, 0, 5684, 23847, 26905, 35080, 15898, 0, 3415, 841, 2677, 2083, 2768, 1774, 1551, 1267, 2045, 482, 3458, 0, 16986, 34892, 28732, 28671, 30241, 16517, 610, 3770, 2003, 3126, 2869, 3224, 3048, 3023, 3175, 3167, 3009, 3009, 3093, 3121, 3030, 3023, 2690, 2471, 2618, 3020, 3459, 3735, 3792, 3816, 3997, 3878, 3994, 4003, 3619, 3463, 1141, 0, 121, 0, 20, 0, 0, 91, 0, 332, 0, 3704, 14398, 18858, 18412, 17662, 17741, 16956, 15843, 15881, 15817, 16063, 14122, 15872, 6710, 0, 812, 0, 208, 43, 967, 1398, 1692, 1812, 1846, 1651, 1433, 1712, 1781, 1968, 2149, 2030, 1145, 814, 421, 0, 57, 0, 15, 0, 1, 0, 0, 9, 0, 33, 0, 313, 999, 1416, 2191, 2634, 2817, 2959, 3049, 3225, 3344, 3453, 3425, 3473, 3632, 3727, 3827, 3936, 4091, 4172, 4059, 4239, 4606, 4849, 5205, 5542, 5732, 5629, 5431, 5072, 3293, 1333, 876, 962, 1021, 968, 1064, 885, 1217, 553, 2739, 5031, 4732, 5125, 4946, 5138, 4968, 4731, 4531, 4331, 4137, 4159, 4071, 3740, 3322, 3359, 3452, 3338, 3381, 3336, 2750, 2084, 1366, 303, 0, 23, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 882, 0, 3133, 0, 20570, 20874, 0, 4112, 0, 1923, 444, 446, 0, 27, 0, 3, 2, 0, 136, 379, 895, 1452, 1589, 1866, 1974, 1747, 1664, 1699, 1648, 1738, 1574, 1898, 838, 0, 100, 0, 17, 4, 0, 330, 1182, 1759, 2236, 2625, 2919, 3001, 2899, 2951, 2668, 2456, 1985, 491, 0, 41, 0, 12, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 32, 0, 111, 0, 972, 2649, 2604, 3054, 2030, 979, 0, 1261, 0, 9133, 24363, 26348, 29583, 30569, 31690, 31781, 31730, 31842, 32005, 31405, 32624, 28309, 27520, 12071, 0, 2461, 463, 1880, 2846, 4012, 3834, 4052, 4100, 3973, 3496, 3373, 3618, 3521, 3582, 3529, 3594, 3485, 3795, 3877, 3573, 3754, 3817, 3829, 3788, 3745, 3737, 3666, 3599, 3573, 3615, 3569, 3567, 3481, 3330, 3210, 3362, 1243, 0, 141, 0, 40, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 28, 0, 332, 1330, 1590, 1584, 1516, 1674, 1336, 2488, 3793, 3550, 3392, 3229, 3524, 3418, 3382, 3413, 3192, 3227, 3258, 3191, 3413, 3492, 3623, 3761, 3737, 3888, 4161, 4142, 4085, 4051, 3836, 3346, 3236, 3076, 2717, 945, 0, 105, 0, 29, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 77, 0, 390, 0, 1373, 0, 11795, 29353, 29610, 33454, 31206, 33521, 30205, 36285, 16797, 0, 3122, 434, 1646, 1409, 0, 2435, 0, 15926, 37344, 27317, 30988, 12299, 0, 2029, 0, 987, 405, 1746, 2263, 2231, 2890, 3308, 3414, 3351, 3456, 3684, 3817, 3770, 3787, 3922, 3710, 3807, 3910, 3830, 3839, 3647, 3527, 3599, 3490, 3682, 3336, 4022, 1778, 0, 221, 0, 63, 0, 12, 0, 40, 0, 194, 0, 673, 0, 6022, 16997, 17617, 18882, 18911, 19249, 19312, 19518, 19550, 19579, 19137, 20055, 18111, 20863, 9000, 0, 1107, 0, 316, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 217, 0, 758, 0, 16596, 30906, 30332, 30577, 34703, 19023, 0, 20098, 32597, 37283, 13143, 11273, 39126, 26060, 33708, 13560, 0, 2862, 725, 2066, 1375, 1986, 2783, 3127, 3339, 3142, 2892, 3031, 2888, 2739, 3035, 3242, 3176, 3226, 3168, 3257, 3090, 3629, 4159, 3873, 3804, 3507, 3070, 2916, 2521, 2311, 871, 0, 101, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 81, 0, 402, 0, 1409, 0, 11718, 28647, 26663, 30020, 30455, 31629, 31355, 31551, 31571, 31066, 30417, 28552, 28396, 26230, 26195, 11232, 0, 1756, 0, 963, 562, 774, 679, 727, 689, 773, 439, 0, 511, 1008, 1023, 966, 1072, 479, 0, 59, 0, 16, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 75, 0, 215, 0, 2868, 13584, 17992, 19553, 7563, 0, 894, 0, 259, 0, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 11, 0, 40, 0, 406, 1395, 1901, 2173, 2171, 2345, 2608, 2593, 1813, 1180, 1314, 1385, 1566, 1981, 2128, 2096, 2112, 2099, 2117, 2087, 2138, 2000, 2008, 755, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 888, 0, 3151, 0, 20634, 20615, 0, 4440, 0, 705, 0, 122, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 110, 0, 378, 0, 4553, 18986, 25749, 27620, 28802, 29193, 30054, 30510, 30473, 30418, 30583, 30316, 30735, 29932, 31430, 28669, 34176, 16076, 0, 3021, 368, 2948, 3010, 3363, 3664, 3756, 3619, 3561, 3509, 3325, 3350, 3447, 3154, 3133, 3014, 3176, 2620, 1945, 789, 0, 109, 0, 107, 66, 0, 9, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 65, 0, 402, 0, 2095, 0, 10066, 22600, 23870, 29521, 29200, 29941, 28968, 30543, 27737, 33306, 14982, 0, 1769, 0, 507, 0, 113, 0, 0, 6, 0, 15, 50, 995, 1928, 2099, 2239, 2358, 2379, 2523, 2592, 2501, 2534, 2592, 2648, 2707, 2826, 2905, 2989, 2970, 2519, 2033, 689, 0, 76, 0, 21, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 24, 0, 186, 548, 1323, 690, 0, 90, 0, 28, 0, 23, 21, 0, 37, 86, 246, 328, 302, 346, 351, 363, 377, 387, 387, 381, 437, 322, 248, 155, 332, 1203, 1815, 1971, 2117, 2233, 2180, 2767, 3194, 3208, 2741, 2347, 2412, 2473, 2275, 2721, 1208, 0, 149, 0, 42, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 29, 0, 102, 0, 867, 2194, 2095, 2289, 2223, 2257, 1934, 1065, 194, 0, 12, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 205, 0, 755, 0, 5693, 11916, 14135, 15007, 10541, 12516, 11093, 9727, 4226, 4515, 3074, 0, 447, 0, 122, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 41, 0, 153, 0, 1751, 7043, 9617, 7551, 6733, 5258, 1676, 2202, 5060, 4626, 10245, 20028, 24065, 26126, 27336, 27901, 27230, 27169, 27967, 29473, 30372, 30442, 30412, 30115, 26670, 24265, 22624, 20176, 17965, 17313, 17526, 18839, 16302, 9558, 8059, 8363, 8064, 8540, 7713, 9320, 4114, 0, 511, 0, 146, 0, 29, 0, 0, 0, 0, 0, 0, 17, 0, 84, 0, 293, 0, 2501, 6711, 6230, 5797, 3481, 4521, 2289, 8909, 16936, 15675, 16388, 16342, 18511, 17837, 18300, 18347, 17557, 13994, 10226, 10441, 10315, 10179, 10642, 9681, 11653, 5156, 0, 640, 0, 183, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 69, 431, 644, 742, 685, 399, 481, 823, 86, 983, 0, 5692, 10953, 9889, 9540, 11287, 7217, 20170, 25583, 12583, 15032, 9033, 7826, 9784, 11127, 12808, 11421, 11264, 10717, 10489, 9175, 7976, 5362, 3698, 3476, 3417, 1622, 0, 178, 0, 48, 0, 9, 0, 0, 0, 0, 0, 7, 0, 36, 0, 127, 0, 987, 2052, 1510, 1793, 1559, 1837, 1391, 2433, 1295, 0, 116, 2078, 5642, 7025, 8007, 9701, 11444, 11634, 11753, 11510, 9752, 8859, 9637, 11475, 14007, 11131, 8123, 6267, 1555, 745, 360, 311, 882, 404, 247, 0, 63, 0, 12, 0, 2, 0, 0, 0, 0, 6, 0, 38, 0, 138, 0, 1319, 4725, 7978, 12775, 13553, 13499, 11502, 3182, 259, 690, 1339, 2796, 1989, 601, 0, 58, 0, 7, 5, 0, 42, 73, 2093, 3873, 4279, 4950, 5702, 6686, 6690, 6430, 5702, 5194, 4512, 4552, 1789, 0, 211, 0, 72, 0, 70, 0, 199, 0, 1658, 4042, 2903, 3247, 2833, 3099, 1413, 0, 182, 0, 50, 0, 10, 0, 3, 0, 12, 0, 97, 46, 47, 0, 256, 0, 1920, 3391, 3963, 6434, 7660, 7128, 10959, 2905, 4302, 6074, 0, 1072, 0, 248, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 68, 0, 246, 0, 2012, 4692, 4317, 4692, 5950, 7098, 6824, 6812, 7082, 6456, 7773, 3418, 0, 368, 284, 1129, 600, 1186, 2003, 1968, 1434, 1828, 792, 0, 96, 0, 28, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 121, 0, 415, 0, 4088, 12890, 12901, 14761, 19810, 21873, 20743, 19588, 19598, 19436, 19393, 19527, 19836, 19377, 18543, 12107, 7801, 11360, 12229, 12830, 12169, 11251, 14111, 14044, 16270, 17449, 15143, 13980, 12505, 9817, 11917, 6140, 0, 653, 0, 182, 0, 35, 0, 0, 0, 0, 0, 3, 0, 39, 0, 170, 0, 884, 312, 4381, 11740, 15297, 24969, 31167, 31132, 29592, 28737, 29857, 30595, 30184, 29970, 30384, 30410, 30526, 30072, 30236, 29910, 29404, 28829, 28807, 27846, 29167, 29884, 28950, 24792, 20323, 20653, 20406, 20385, 20747, 19882, 21637, 17306, 18249, 7989, 7452, 21938, 6470, 0, 553, 0, 197, 0, 55, 0, 0, 0, 1, 0, 8, 0, 96, 301, 985, 650, 906, 46, 3275, 6333, 6277, 3531, 0, 223, 0, 62, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 15, 155, 0, 393, 0, 1133, 0, 8176, 15898, 7603, 5346, 0, 4703, 16100, 6850, 0, 681, 0, 211, 0, 50, 0, 4, 0, 8, 61, 961, 2277, 2539, 2984, 1753, 569, 1179, 966, 1363, 629, 0, 80, 0, 23, 0, 4, 0, 0, 0, 12, 0, 62, 0, 247, 0, 1855, 3431, 3457, 1619, 6148, 17726, 22214, 22503, 23612, 26116, 27201, 29063, 30286, 30380, 29973, 29970, 29709, 29324, 28694, 28019, 28400, 27963, 28080, 27879, 27810, 23936, 19327, 18637, 16668, 16442, 16388, 13997, 13873, 14585, 14853, 13400, 13850, 5619, 0, 674, 0, 192, 0, 38, 0, 0, 0, 0, 0, 0, 2, 0, 5, 0, 78, 291, 120, 69, 300, 506, 931, 1379, 2318, 2503, 2760, 2911, 2416, 2244, 1502, 594, 5, 140, 529, 833, 3837, 6364, 4259, 3199, 4159, 5286, 5516, 4585, 4330, 4419, 4286, 4523, 4096, 4939, 2183, 0, 271, 0, 77, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 25, 0, 92, 0, 744, 1672, 1476, 1719, 2073, 1799, 1276, 1370, 1353, 1237, 1239, 704, 422, 290, 0, 43, 0, 11, 0, 1, 0, 0, 0, 1, 0, 11, 0, 47, 0, 289, 403, 1390, 2558, 2599, 2780, 2785, 2774, 3054, 3889, 3421, 939, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 5, 0, 8, 188, 2250, 4278, 4425, 4475, 4407, 4507, 4338, 4669, 3597, 2534, 2563, 2355, 2193, 1826, 1836, 1368, 671, 383, 237, 0, 11, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 232, 0, 826, 0, 5958, 10633, 10866, 19640, 17630, 15771, 16922, 16719, 17384, 16932, 18171, 23117, 25817, 27413, 26137, 25272, 26110, 26178, 25719, 25425, 26012, 26571, 25891, 24717, 24472, 23396, 22705, 18830, 16639, 13468, 7203, 3726, 1611, 1190, 283, 0, 14, 0, 4, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 9, 0, 0, 0, 500, 3264, 988, 9958, 19170, 17736, 19667, 20324, 21550, 21960, 22013, 22829, 25653, 27297, 27832, 28083, 28581, 28584, 28341, 28033, 27529, 27265, 26931, 27258, 26682, 27755, 25765, 29725, 17239, 7251, 9161, 6124, 3674, 0, 470, 0, 0, 275, 0, 2238, 2461, 0, 330, 0, 182, 0, 647, 627, 0, 95, 0, 30, 0, 41, 0, 869, 2128, 5127, 6526, 11142, 18333, 19668, 21720, 22282, 21067, 22577, 24587, 24961, 25005, 24807, 25207, 24392, 26999, 29269, 28986, 29815, 29855, 30637, 30600, 31331, 31486, 31829, 31793, 31556, 30976, 30895, 30053, 31891, 29651, 34657, 18222, 0, 18966, 33885, 26537, 14672, 1440, 0, 9346, 17965, 16621, 18130, 17377, 17612, 17484, 15178, 17989, 7468, 0, 0, 5168, 12642, 9993, 11610, 10246, 12017, 6624, 0, 2232, 271, 12169, 25652, 25330, 29120, 28048, 29250, 17774, 8247, 11341, 9906, 10665, 8625, 8048, 5635, 2054, 784, 0, 96, 0, 21, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 51, 0, 104, 36, 4107, 10319, 6563, 6571, 1801, 6364, 17267, 18298, 22387, 25284, 28428, 28282, 28589, 29367, 26752, 23107, 19468, 16400, 11406, 6390, 6131, 5137, 3479, 2787, 3152, 2898, 2476, 1662, 1355, 1443, 1371, 1464, 1318, 1594, 703, 0, 87, 0, 25, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 89, 0, 315, 0, 2588, 6239, 6334, 8242, 8723, 5358, 2485, 1525, 8491, 18328, 20552, 25313, 27401, 25646, 26323, 24111, 22094, 22938, 22043, 23368, 21114, 25488, 11267, 0, 1400, 0, 400, 0, 81, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 31, 0, 100, 0, 1073, 4269, 5578, 7728, 7459, 15349, 20913, 18814, 19097, 18115, 17326, 20077, 24507, 24551, 24656, 24721, 24448, 25024, 23845, 27964, 33250, 31669, 32704, 29321, 24101, 23580, 13485, 6417, 6908, 5110, 4733, 3102, 2233, 1874, 623, 0, 65, 0, 18, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 73, 0, 357, 0, 1243, 0, 9917, 21466, 14752, 13655, 11834, 10876, 9371, 8372, 7412, 5216, 3411, 4153, 3780, 4050, 2629, 6717, 9739, 10489, 8005, 4429, 5039, 4015, 3236, 1602, 564, 0, 45, 0, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 152, 0, 543, 0, 5670, 9981, 9283, 10230, 8385, 9787, 10515, 11115, 10611, 10558, 10299, 8646, 6695, 5931, 3780, 11148, 20766, 22641, 24809, 25909, 26939, 27274, 28407, 29827, 30150, 30674, 30087, 30105, 25526, 22023, 19983, 19499, 14199, 7374, 7435, 6004, 5152, 4411, 4690, 4469, 4752, 4293, 5184, 2291, 0, 284, 0, 81, 0, 16, 0, 0, 0, 0, 0, 0, 2, 0, 13, 0, 67, 0, 522, 1043, 1891, 956, 4577, 8732, 7824, 10094, 10448, 15118, 18485, 17515, 17090, 15468, 13193, 11189, 11400, 11383, 10040, 9045, 9372, 9138, 9402, 9006, 9743, 7404, 4996, 4609, 3634, 3846, 3262, 3184, 3270, 3886, 1469, 0, 168, 0, 48, 0, 10, 0, 0, 0, 0, 18, 0, 80, 0, 269, 0, 3192, 12623, 15090, 16581, 20683, 23358, 24555, 25075, 26382, 27437, 27288, 25299, 24343, 24635, 24399, 24696, 24230, 25100, 22343, 20069, 21952, 21292, 21955, 21643, 20393, 20703, 21485, 21642, 21301, 21006, 19454, 17807, 13675, 11448, 11299, 11707, 11835, 11049, 4095, 0, 470, 0, 133, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 0, 183, 0, 641, 0, 4491, 6113, 0, 438, 0, 151, 20, 561, 2335, 5224, 7086, 8128, 8411, 8252, 9031, 9381, 8216, 8021, 2911, 0, 330, 0, 95, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 118, 0, 419, 0, 3717, 10608, 12477, 14923, 15023, 15282, 14118, 15917, 11995, 12404, 20053, 23756, 27030, 27008, 27731, 25951, 19880, 12877, 13441, 5641, 0, 682, 0, 194, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 19, 113, 28, 332, 769, 2583, 3224, 4497, 9641, 10800, 10847, 12862, 12810, 17825, 22041, 20939, 20315, 18611, 17896, 18270, 17707, 18687, 16923, 20406, 9025, 0, 1121, 0, 320, 0, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 178, 0, 667, 0, 5217, 12455, 18295, 22394, 19505, 20617, 19101, 16458, 4923, 0, 492, 0, 14, 47, 1701, 15787, 9224, 0, 1750, 1683, 3268, 4237, 6799, 5268, 1597, 0, 267, 0, 82, 0, 16, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 9, 0, 7, 0, 291, 1841, 450, 439, 0, 4977, 11977, 13695, 19168, 23379, 27581, 28586, 29640, 29627, 27597, 26364, 24339, 25232, 18014, 9775, 3919, 0, 506, 0, 131, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 117, 0, 415, 0, 3628, 7634, 7771, 11419, 12552, 11660, 9666, 4698, 563, 608, 699, 855, 1293, 1954, 1968, 986, 706, 1749, 1845, 3169, 7802, 9855, 9090, 8509, 6933, 6718, 6701, 6394, 6299, 5809, 5779, 5638, 5928, 5382, 6481, 2869, 0, 356, 0, 101, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 141, 0, 523, 0, 4217, 10530, 15465, 19414, 19007, 18728, 21580, 6869, 4134, 20548, 22535, 25924, 26835, 28401, 28513, 28207, 28729, 28814, 29128, 28373, 29853, 27085, 32629, 14438, 0, 1793, 0, 513, 0, 104, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 105, 0, 450, 0, 1539, 0, 12264, 28172, 25421, 29046, 26537, 26787, 22736, 21784, 18375, 14959, 6466, 0, 656, 0, 180, 0, 32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 13, 0, 104, 0, 1211, 660, 1889, 0, 8500, 13572, 15123, 8738, 0, 1445, 1834, 6217, 7720, 9123, 7994, 6985, 7011, 6624, 7044, 6258, 6531, 3502, 0, 158, 0, 48, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 335, 4507, 13534, 17441, 16649, 16754, 15511, 14626, 14166, 13585, 12586, 11851, 10862, 9562, 5748, 2746, 4606, 5911, 6500, 7671, 8452, 9078, 8796, 8307, 7782, 7189, 7094, 6621, 6607, 6825, 6850, 6929, 6746, 7101, 6442, 7761, 3434, 0, 426, 0, 122, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16370, 11030, 12858, 15138, 23738, 18804, 13682, 9800, 13808, 7272, 13468, 7074, 6450, 12008, 2710, 5132, 13168, 13118, 16014, 19942, 31802, 15382, 0, 10594, 24200, 28806, 30646, 32186, 32502, 32252, 33182, 33008, 32784, 33424, 32136, 34788, 25428, 13094, 17536, 15026, 21010, 33112, 28030, 22386, 24806, 24166, 23190, 24710, 27986, 27788, 34234, 32764, 29856, 14564, 0, 11816, 22546, 22820, 26944, 27522, 30826, 26422, 28064, 27760, 28638, 26704, 25782, 23884, 3860, 686, 72, 2914, 7622, 15288, 22218, 20142, 21040, 20800, 20504, 21616, 16416, 3534, 0, 802, 0, 3950, 5454, 7304, 8512, 4290, 2384, 0, 364, 0, 192, 0, 402, 0, 2608, 2428, 0, 0, 750, 0, 6240, 6394, 0, 1216, 0, 1466, 0, 3474, 3700, 0, 578, 0, 160, 0, 22, 12, 0, 76, 0, 224, 0, 2188, 4848, 0, 7286, 23448, 22588, 27654, 20560, 17266, 21248, 10700, 16558, 10586, 0, 11626, 7250, 6824, 4926, 5948, 8948, 378, 15708, 5002, 294, 7532, 10680, 10056, 3708, 8158, 16548, 17798, 16782, 19558, 22180, 27244, 31936, 32946, 34990, 34602, 34148, 35570, 32662, 38626, 18648, 0, 1982, 0, 2058, 1470, 0, 994, 658, 0, 132, 0, 246, 0, 756, 0, 6030, 10004, 2902, 1022, 0, 0, 1430, 1150, 434, 1438, 0, 1194, 0, 5582, 2170, 5944, 7762, 0, 774, 260, 0, 7490, 17216, 14442, 15428, 15600, 14210, 17832, 8070, 0, 422, 2534, 11182, 6254, 246, 134, 0, 116, 0, 68, 0, 266, 0, 3094, 13156, 22986, 27308, 28796, 30898, 30856, 31470, 31700, 32052, 30850, 26972, 19538, 14538, 8554, 5028, 6642, 5962, 6556, 6324, 5280, 5022, 5562, 5610, 5772, 5442, 6058, 4750, 10130, 23218, 29496, 32106, 35036, 35560, 35448, 33626, 32638, 33636, 24602, 23362, 34246, 19526, 4950, 6936, 5888, 8346, 6846, 5472, 7140, 5106, 5156, 4702, 1132, 3142, 4410, 5380, 4684, 13260, 14968, 11752, 17988, 16538, 18512, 21430, 10900, 456, 212, 0, 228, 0, 562, 0, 3444, 3002, 1566, 15196, 19652, 25920, 29526, 26868, 35438, 26824, 17502, 14170, 8216, 15836, 6302, 0, 928, 756, 2080, 3164, 11334, 14198, 15336, 12742, 8256, 5028, 860, 0, 1434, 9914, 15028, 14964, 15432, 6288, 7570, 20656, 25730, 28636, 30332, 30366, 30502, 30308, 30610, 30018, 32124, 34298, 28120, 18172, 15986, 16328, 22830, 29840, 26124, 25658, 31512, 30522, 24222, 25256, 30006, 32396, 33716, 27964, 32558, 11054, 5628, 24388, 18662, 24784, 25776, 28768, 33452, 33868, 24808, 25988, 31762, 32628, 23142, 24524, 20018, 4324, 17198, 8188, 0, 1018, 0, 342, 0, 138, 0, 3238, 21718, 27102, 6682, 0, 336, 38, 0, 4380, 3806, 0, 0, 802, 0, 6652, 7416, 0, 2698, 0, 11062, 10606, 0, 1744, 0, 1348, 0, 4978, 0, 24938, 11432, 20434, 19960, 12542, 25880, 0, 4860, 0, 1012, 0, 304, 0, 586, 0, 5014, 13644, 18164, 17054, 12092, 12682, 17378, 16080, 24692, 29132, 0, 16326, 18068, 518, 0, 15996, 14992, 32, 7372, 0, 14438, 4130, 11188, 25954, 27994, 21528, 20532, 17344, 13760, 21690, 22212, 23972, 20544, 20760, 21966, 25950, 28930, 29170, 29250, 29510, 28802, 30232, 27544, 32934, 15152, 0, 1744, 0, 764, 0, 1856, 1348, 290, 1204, 0, 738, 0, 2922, 1308, 12160, 10922, 5852, 6474, 0, 1070, 0, 270, 0, 12, 54, 0, 300, 0, 1460, 0, 3734, 3972, 0, 234, 396, 0, 5896, 13460, 11280, 12114, 12114, 11290, 13426, 5978, 0, 740, 0, 210, 0, 42, 0, 0, 0, 14, 0, 90, 0, 1682, 10314, 22106, 27000, 31474, 35908, 35256, 35458, 34866, 36226, 34718, 34098, 26210, 24868, 24358, 15724, 10298, 6214, 7852, 6594, 6702, 4964, 4476, 5580, 5452, 5274, 5908, 4572, 7108, 2004, 19010, 37834, 34136, 36804, 34214, 34160, 34560, 29398, 32804, 21558, 22232, 32266, 14190, 7112, 5612, 8884, 9522, 6766, 7832, 7328, 6606, 6892, 5660, 4996, 6306, 4466, 5528, 7054, 18560, 18000, 13604, 17670, 17876, 17776, 10086, 5210, 1580, 0, 10, 26, 0, 312, 0, 1190, 0, 9822, 24004, 28182, 29054, 31570, 30874, 31030, 28152, 26330, 16666, 11368, 16778, 4922, 0, 12206, 21296, 15130, 18854, 16448, 19868, 18186, 18590, 4624, 3978, 12200, 5582, 10074, 12564, 17206, 14638, 12986, 4072, 5826, 22188, 25692, 30952, 31092, 31050, 31056, 31024, 31066, 31022, 31092, 30838, 30696, 30900, 32542, 30166, 34614, 31138, 24294, 25232, 22092, 20232, 17224, 21054, 24002, 28090, 30414, 33166, 14602, 1116, 3964, 2408, 3228, 16786, 31796, 34226, 36570, 34770, 32374, 31012, 29136, 27418, 27244, 22990, 32946, 11866, 8752, 11236, 0, 1870, 0, 470, 0, 0, 462, 0, 1752, 0, 12642, 11808, 0, 910, 2682, 11658, 16158, 7280, 0, 1304, 0, 1782, 0, 10068, 10666, 0, 3050, 0, 10510, 12438, 0, 11586, 2330, 10500, 4258, 14734, 14140, 7408, 19572, 0, 17268, 12742, 0, 1842, 0, 574, 0, 74, 38, 0, 144, 814, 11458, 14764, 0, 7810, 21438, 25838, 25920, 24534, 19826, 26768, 23678, 25556, 21214, 3006, 0, 13140, 12914, 0, 3196, 25636, 18084, 0, 2936, 0, 2362, 0, 10850, 26354, 23882, 26162, 28210, 28492, 24536, 24162, 22404, 29400, 31374, 26864, 29000, 26938, 29868, 24910, 34248, 8968, 13238, 20974, 0, 330, 5614, 8698, 0, 8, 3066, 3484, 0, 0, 1256, 0, 12316, 25090, 6230, 652, 0, 1182, 0, 8452, 16272, 21612, 22370, 3890, 0, 1466, 0, 9394, 10986, 0, 7316, 0, 11060, 12268, 0, 2112, 0, 1352, 0, 2970, 0, 18874, 18702, 0, 2416, 0, 0, 5234, 6850, 0, 5506, 3646, 0, 0, 3160, 4008, 10288, 21474, 25070, 30992, 34510, 37310, 36860, 35442, 33136, 34524, 34106, 23582, 16304, 17796, 25408, 31584, 23506, 9466, 8792, 4010, 17646, 16482, 6734, 16026, 11952, 14460, 12466, 14748, 10942, 23178, 37988, 37708, 40752, 39724, 38642, 38982, 37686, 34702, 34388, 34588, 30368, 31422, 20724, 12392, 27216, 22386, 10918, 8358, 7126, 6550, 6360, 5952, 5520, 2798, 9188, 15368, 22754, 14442, 0, 6196, 18368, 19810, 17826, 19350, 14108, 2844, 1788, 5998, 4510, 5362, 4664, 5512, 4186, 6256, 0, 10012, 20698, 22876, 32688, 32332, 27074, 20432, 23952, 16634, 3084, 0, 518, 0, 252, 0, 602, 0, 9896, 12470, 13382, 9668, 266, 0, 3124, 1894, 4554, 17376, 16018, 21194, 16114, 12820, 2026, 11026, 31238, 32578, 36254, 33626, 34798, 34172, 34586, 34168, 34836, 33084, 32812, 30188, 31410, 34446, 33386, 26478, 26606, 26830, 21728, 23872, 21742, 23080, 24718, 25776, 27016, 35226, 15754, 0, 5812, 0, 12884, 29722, 32046, 38376, 32374, 33588, 23706, 28724, 16104, 17916, 27662, 27692, 14066, 17440, 12890, 8474, 18690, 0, 6466, 0, 6614, 0, 22726, 20582, 0, 2600, 0, 0, 6902, 14520, 19886, 28750, 28320, 10734, 0, 162, 1422, 0, 12482, 10014, 3202, 12928, 0, 18394, 8856, 11032, 16940, 0, 2990, 0, 1348, 0, 2208, 0, 13664, 13648, 0, 2042, 0, 408, 364, 1464, 1236, 1096, 1558, 500, 4968, 16334, 20786, 20800, 14976, 22044, 27134, 30670, 28638, 29074, 24688, 24100, 29862, 28328, 6620, 10614, 18544, 0, 20120, 18548, 0, 11768, 4490, 5698, 8032, 0, 742, 1006, 320, 4906, 17576, 22122, 23758, 27474, 28474, 23374, 24278, 24346, 24008, 24968, 23836, 25770, 22278, 29022, 9666, 5308, 10020, 0, 1732, 0, 528, 0, 458, 0, 1420, 0, 9196, 8824, 0, 468, 3858, 15890, 5764, 0, 170, 1612, 6538, 10630, 15164, 6532, 0, 3648, 0, 19922, 20290, 0, 4612, 0, 11274, 10008, 0, 1538, 0, 432, 0, 24, 92, 0, 428, 0, 4022, 12558, 13928, 4912, 0, 562, 0, 278, 0, 524, 0, 3402, 6302, 13318, 21662, 24558, 30844, 31510, 33238, 34124, 33100, 32750, 32966, 30470, 27350, 25734, 29362, 16938, 5228, 7756, 6410, 7234, 6502, 6866, 4422, 8922, 13696, 12012, 13276, 11834, 13998, 9988, 22828, 35864, 33986, 38280, 35708, 35730, 35244, 31592, 27582, 28182, 25526, 15654, 8204, 6274, 6588, 6840, 6408, 6546, 6754, 7110, 3770, 3122, 5312, 6380, 4354, 9378, 10490, 14918, 11066, 0, 16192, 22936, 13696, 5858, 0, 9802, 9684, 1390, 0, 48, 0, 306, 0, 1088, 0, 9598, 26364, 27162, 25844, 26400, 24756, 23900, 30674, 18074, 6482, 2758, 0, 464, 0, 810, 0, 3938, 8616, 15778, 16986, 20988, 11470, 0, 12726, 2560, 5858, 18492, 14918, 21436, 15870, 13122, 2994, 9166, 30496, 31106, 33366, 32008, 32832, 32480, 32636, 32574, 32594, 32608, 32348, 30874, 30252, 35154, 31714, 26146, 27538, 24718, 24096, 23790, 22682, 24414, 27708, 27274, 33902, 13376, 0, 9434, 3768, 0, 10328, 27616, 30442, 35734, 33738, 31990, 26452, 28120, 22856, 30240, 14528, 15792, 20166, 10692, 8518, 2690, 10700, 424, 2562, 1296, 1702, 2026, 864, 3198, 0, 19096, 13940, 0, 148, 6222, 18042, 23574, 30242, 28548, 10074, 0, 0, 4686, 5120, 0, 3836, 0, 6466, 6516, 0, 3356, 0, 11802, 6268, 8768, 12940, 0, 1394, 2102, 0, 18316, 18052, 0, 2722, 0, 768, 0, 230, 0, 398, 0, 1476, 0, 11344, 22222, 16184, 3270, 8464, 23936, 23136, 15368, 17756, 13886, 24136, 17120, 0, 1052, 7056, 32428, 16550, 21900, 18826, 0, 650, 956, 0, 12470, 17416, 15164, 32780, 20968, 19862, 24630, 25706, 23466, 23970, 28656, 24586, 21432, 20814, 19366, 18350, 18832, 18214, 19240, 17416, 21008, 9290, 0, 1154, 0, 330, 0, 66, 0, 34, 0, 186, 0, 660, 0, 4320, 4350, 0, 772, 0, 532, 0, 3158, 10056, 13394, 20658, 9194, 0, 2456, 0, 13146, 32646, 9272, 0, 3238, 0, 2502, 0, 15806, 35022, 29664, 31470, 32114, 28840, 36366, 13066, 7382, 31450, 2942, 9830, 11630, 0, 5840, 4098, 0, 5338, 8084, 5604, 11270, 11774, 15108, 21640, 26342, 29682, 31004, 32158, 32106, 31406, 29794, 29640, 25228, 19590, 21716, 14314, 6230, 7160, 5936, 7576, 5018, 11666, 9746, 2446, 5286, 3858, 4336, 4606, 3496, 5834, 1020, 17070, 34760, 32364, 36494, 35966, 36738, 35500, 33444, 33308, 34554, 25780, 24550, 18698, 5910, 8336, 9074, 7268, 6956, 6640, 7312, 4696, 3966, 3940, 1840, 3166, 2992, 3942, 0, 10754, 4682, 10696, 23214, 12750, 11200, 0, 9284, 7138, 0, 1010, 0, 118, 194, 0, 1182, 0, 10464, 26598, 20038, 20030, 23194, 21114, 22406, 18782, 9954, 15902, 13320, 7970, 11696, 9090, 0, 11792, 21036, 15132, 16822, 9812, 22514, 22166, 20280, 24988, 18098, 17362, 19840, 20120, 20740, 15900, 5286, 0, 11022, 26556, 26006, 27592, 30866, 34364, 33594, 33314, 34690, 31700, 37716, 20600, 20232, 30122, 18296, 26394, 29658, 34962, 24722, 18502, 22904, 19260, 18898, 21010, 24152, 32580, 13148, 0, 2006, 0, 1744, 0, 10832, 27810, 29608, 31564, 27284, 29462, 28254, 27494, 35350, 23046, 17340, 20754, 10950, 0, 16204, 17078, 6458, 18216, 13574, 15692, 15160, 14344, 16976, 7552, 0, 894, 0, 108, 94, 464, 9730, 14484, 3458, 0, 220, 0, 0, 318, 0, 1256, 0, 8516, 9358, 0, 4928, 2858, 0, 452, 0, 582, 0, 1608, 0, 10480, 10650, 0, 2086, 480, 6298, 28000, 14968, 0, 1712, 0, 0, 1172, 0, 11226, 20632, 6454, 0, 9342, 15436, 6856, 7732, 3216, 5836, 6058, 0, 14026, 12168, 0, 0, 6824, 8414, 0, 1074, 0, 0, 1850, 0, 24152, 20950, 15692, 19064, 13792, 27568, 20124, 24630, 19384, 16190, 20556, 19974, 20806, 12570, 4556, 7086, 5688, 6674, 5730, 7090, 3096, 0, 408, 0, 176, 0, 26, 20, 1078, 5792, 0, 20488, 19820, 0, 2836, 0, 282, 602, 0, 8076, 18982, 15084, 31280, 16924, 0, 2438, 0, 13820, 12122, 0, 11346, 9338, 0, 2358, 0, 5644, 0, 14646, 36140, 28648, 33386, 29266, 34578, 18728, 0, 5692, 0, 26524, 17782, 12418, 34846, 6182, 21422, 15426, 10852, 9820, 11330, 8254, 0, 11912, 24916, 25100, 29180, 28758, 28706, 26466, 27000, 27534, 27650, 23284, 30948, 21288, 7734, 8558, 9524, 19160, 12090, 4916, 3362, 6224, 7056, 9114, 12890, 11988, 11820, 13034, 10086, 20196, 30874, 31410, 35262, 33750, 34354, 32440, 30834, 32998, 29190, 27150, 19140, 15370, 11108, 13212, 11050, 3638, 7452, 3092, 4694, 1226, 744, 2168, 0, 4532, 4098, 0, 2092, 0, 8942, 4616, 8954, 25880, 1998, 6502, 6098, 0, 0, 6250, 15642, 12870, 13708, 14226, 12228, 17084, 6652, 4244, 21332, 8270, 12786, 17772, 19678, 21832, 18290, 5998, 3706, 9292, 0, 13896, 20658, 6424, 15802, 21680, 21564, 22504, 24552, 23234, 17052, 17038, 19922, 21826, 25126, 25622, 16620, 4996, 0, 8456, 21008, 21480, 23460, 23604, 27580, 29446, 29026, 29118, 29304, 28732, 29950, 26778, 27904, 24508, 19454, 23086, 18694, 17062, 17176, 17682, 17068, 17452, 14008, 2670, 0, 0, 2160, 2882, 0, 1662, 0, 10604, 25490, 23252, 24206, 24476, 26712, 15492, 20962, 23658, 24640, 26358, 18138, 7386, 0, 916, 0, 238, 0, 42, 0, 0, 0, 76, 0, 402, 0, 1404, 0, 15676, 33938, 32282, 31390, 25294, 9326, 0, 2160, 720, 0, 734, 0, 2732, 0, 16212, 10604, 7852, 14414, 0, 2482, 0, 588, 0, 0, 740, 0, 2568, 0, 18754, 31222, 4562, 19676, 5608, 19338, 44428, 36412, 40082, 38906, 37962, 41748, 27212, 7434, 2130, 2944, 14770, 23244, 11926, 17644, 10838, 17380, 3404, 20984, 17692, 12082, 26242, 0, 30912, 35260, 38262, 28056, 30458, 35942, 42544, 25356, 14990, 43398, 21812, 23364, 25048, 21102, 20266, 17256, 16552, 16540, 17432, 9714, 7174, 13714, 13746, 14382, 13456, 15058, 12126, 17740, 3232, 10520, 13520, 0, 3302, 0, 4922, 0, 25096, 25190, 0, 3856, 0, 1054, 0, 98, 120, 0, 954, 946, 5170, 18110, 7882, 0, 220, 848, 0, 8836, 9236, 0, 2102, 0, 2962, 0, 16944, 16944, 9244, 8186, 9335, 8675, 8601, 6693, 4002, 1908, 1181, 1682, 2332, 2993, 3451, 4618, 4460, 4401, 4101, 4817, 3404, 6053, 704, 18440, 35106, 18992, 4920, 7867, 17969, 18981, 18912, 18526, 20964, 20809, 21043, 20554, 20642, 20131, 20774, 18267, 15116, 16549, 17642, 17867, 18249, 18559, 17529, 17951, 18092, 17910, 18127, 18300, 13993, 5844, 6313, 3520, 0, 334, 0, 97, 0, 25, 0, 45, 0, 190, 0, 1514, 3587, 6398, 8898, 13724, 15829, 14613, 17365, 17225, 18080, 17517, 17920, 14312, 12606, 15405, 9369, 6888, 10118, 2836, 1156, 2434, 0, 1487, 1143, 0, 59, 0, 27, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 35, 0, 112, 0, 1039, 3486, 4672, 7452, 4371, 649, 191, 2695, 6827, 7519, 8991, 9650, 7060, 5098, 5754, 5522, 5525, 5921, 5500, 5864, 7993, 8706, 9606, 10194, 10290, 8468, 8229, 9636, 8014, 9499, 3455, 0, 1279, 0, 257, 0, 62, 0, 35, 0, 139, 0, 486, 0, 4047, 9867, 9027, 10139, 10222, 10431, 10341, 10997, 11134, 11125, 11148, 10934, 11512, 10374, 10294, 11049, 11437, 12413, 13073, 10527, 12185, 5634, 0, 715, 0, 203, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 106, 0, 370, 0, 3189, 8416, 7963, 7878, 7174, 7509, 6824, 6049, 6319, 6569, 6438, 6365, 6624, 6485, 6744, 6855, 6687, 6738, 7016, 7000, 7488, 7430, 6296, 5782, 6609, 7140, 8854, 3700, 0, 444, 0, 149, 0, 138, 0, 382, 0, 4950, 9745, 8411, 8896, 8963, 8307, 9948, 4343, 0, 854, 4378, 5109, 2821, 5717, 2132, 0, 236, 0, 76, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 67, 0, 234, 0, 1953, 2255, 0, 182, 0, 53, 0, 7, 0, 22, 0, 132, 0, 454, 0, 5582, 8793, 5459, 6682, 6062, 6140, 5765, 5374, 5543, 5165, 7078, 8495, 10036, 6305, 172, 171, 0, 54, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 23, 0, 73, 0, 785, 2521, 2002, 3997, 6426, 5877, 6635, 7494, 7159, 8217, 3030, 2822, 6182, 7398, 5141, 5314, 3739, 0, 545, 0, 148, 0, 26, 0, 0, 0, 0, 0, 0, 0, 12, 0, 57, 0, 198, 0, 1926, 6173, 6719, 6796, 6602, 6935, 6343, 7521, 3495, 0, 799, 0, 4481, 15728, 11113, 8082, 4276, 0, 607, 0, 169, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 55, 0, 227, 596, 5332, 5688, 1873, 3814, 1314, 475, 1478, 1, 80, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 162, 0, 563, 0, 5070, 14336, 14396, 14913, 15919, 16620, 16523, 16370, 16805, 15922, 17713, 12000, 7046, 7754, 8710, 10887, 8528, 9678, 8960, 7328, 7918, 4871, 1782, 1779, 1294, 1239, 628, 27, 5, 9, 27, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 20, 0, 72, 0, 635, 1783, 2487, 5083, 6818, 6534, 6266, 4630, 4002, 1644, 0, 203, 0, 56, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 22, 369, 5107, 11661, 13183, 13125, 13037, 13874, 13852, 13058, 13306, 13235, 13163, 13409, 12689, 12431, 9093, 2949, 442, 0, 32, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 89, 615, 338, 0, 43, 0, 12, 0, 2, 0, 0, 0, 0, 1, 0, 8, 0, 30, 0, 200, 200, 0, 30, 0, 8, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 21, 0, 106, 0, 1068, 3801, 6545, 1511, 2650, 8278, 9352, 4258, 0, 539, 0, 146, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 170, 0, 601, 0, 4919, 11509, 10652, 10814, 10942, 11454, 13469, 5776, 0, 703, 0, 200, 0, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 161, 0, 563, 0, 4632, 11084, 10119, 11793, 11667, 11504, 11115, 11300, 11446, 11813, 12197, 12622, 13791, 9253, 5936, 6954, 6314, 6907, 6138, 7472, 3288, 0, 409, 0, 117, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 71, 0, 310, 0, 1582, 0, 3699, 6280, 6550, 10694, 9233, 9227, 9001, 9357, 9213, 8681, 8379, 3220, 0, 377, 0, 106, 0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 8, 0, 40, 0, 336, 793, 905, 41, 1619, 2550, 347, 0, 0, 1, 2, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 28, 0, 102, 0, 1056, 3960, 5727, 5725, 4245, 3572, 3955, 4469, 5436, 5586, 6404, 6946, 7505, 7287, 8128, 3535, 0, 436, 0, 124, 0, 24, 84, 839, 1097, 1001, 461, 0, 53, 0, 35, 0, 184, 490, 754, 852, 908, 820, 1055, 424, 2287, 5276, 5553, 4998, 4863, 4799, 1384, 0, 133, 0, 39, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 32, 0, 85, 0, 1307, 5464, 2490, 0, 298, 0, 90, 0, 20, 0, 0, 0, 0, 0, 0, 0, 8, 0, 50, 0, 189, 0, 1719, 5428, 8932, 12752, 15017, 15325, 14688, 14848, 15329, 15061, 9033, 11384, 5827, 8696, 11153, 3653, 6480, 5005, 5810, 5356, 5683, 5052, 4310, 4797, 4377, 4320, 4235, 5421, 2432, 0, 301, 0, 90, 0, 48, 0, 103, 0, 2123, 2307, 755, 308, 86, 0, 2051, 6093, 6570, 6545, 5875, 5652, 5933, 5663, 6797, 7496, 7278, 7410, 7545, 7489, 6460, 6335, 6402, 6229, 6585, 5910, 7254, 3085, 376, 2115, 1675, 1150, 0, 165, 0, 37, 0, 12, 0, 47, 0, 159, 0, 3273, 2653, 1241, 6827, 9421, 10422, 10214, 9778, 10314, 9079, 6690, 7048, 8686, 8829, 9954, 11547, 11511, 11382, 8786, 8535, 10749, 9307, 8640, 8823, 8650, 8893, 8497, 9275, 6378, 870, 0, 8, 0, 4, 0, 0, 0, 0, 25, 0, 70, 146, 4045, 9178, 9271, 8195, 8568, 8257, 5474, 4815, 6430, 6559, 7105, 7711, 7379, 7420, 6789, 8130, 8289, 8029, 9702, 8126, 9126, 3827, 0, 469, 0, 135, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 166, 1595, 4954, 9690, 10305, 9857, 9303, 10363, 10582, 10158, 13475, 12714, 11897, 12418, 12689, 13190, 13610, 11097, 12299, 9860, 10872, 8628, 2681, 4670, 3590, 4116, 3761, 4076, 3659, 4421, 1956, 0, 253, 0, 111, 0, 135, 0, 1339, 4511, 2964, 6845, 10347, 10477, 11327, 10312, 10159, 12500, 12630, 13828, 9842, 7435, 9861, 8135, 9052, 8700, 9062, 8371, 8743, 9260, 10383, 10011, 9120, 8940, 6408, 8801, 4144, 0, 526, 0, 152, 0, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 55, 0, 197, 0, 2190, 8820, 13341, 15179, 14536, 14184, 14262, 14567, 16343, 14673, 16090, 11352, 11058, 5000, 4434, 5664, 0, 926, 0, 242, 0, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 116, 0, 413, 0, 3459, 8887, 9927, 11254, 10420, 10479, 10305, 10860, 11072, 11450, 11835, 12004, 12292, 12293, 12335, 12167, 12075, 12456, 12419, 11104, 5906, 734, 0, 6, 0, 0, 0, 0, 0, 0, 17, 0, 59, 0, 176, 0, 1928, 5746, 1071, 2570, 10579, 13695, 16357, 18072, 17584, 17044, 18043, 18410, 18348, 19067, 18619, 18874, 16257, 13191, 13220, 13379, 13584, 13516, 12662, 12049, 8771, 10699, 8607, 496, 168, 0, 55, 0, 0, 0, 0, 8, 0, 37, 0, 127, 0, 1599, 6865, 9443, 10527, 11593, 11211, 11569, 12069, 13102, 14067, 11882, 7624, 6480, 6470, 6386, 7152, 6794, 6272, 7133, 6941, 8741, 11810, 12013, 12294, 12558, 12917, 13031, 11730, 8533, 8488, 10185, 11370, 9011, 2083, 0, 163, 0, 50, 0, 11, 0, 0, 0, 0, 0, 0, 8, 0, 52, 0, 206, 0, 2016, 7450, 12741, 13393, 11909, 14262, 11985, 7032, 637, 2135, 2507, 0, 394, 0, 107, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 56, 0, 196, 0, 2103, 7666, 9477, 9594, 10207, 10293, 10290, 10270, 10082, 10046, 7213, 4882, 2053, 0, 1924, 5106, 5611, 5662, 5797, 5898, 6611, 5815, 8878, 11760, 11152, 11641, 11423, 10541, 8376, 9674, 3969, 0, 474, 0, 137, 0, 49, 0, 106, 0, 376, 0, 2859, 5580, 4538, 7219, 8156, 8055, 7807, 7983, 8145, 8600, 8473, 8767, 8729, 8682, 7332, 9178, 3299, 1444, 7660, 8179, 7186, 1527, 0, 113, 0, 41, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 299, 2570, 3862, 3468, 3745, 3441, 3889, 3071, 5589, 7727, 7973, 9777, 9633, 9026, 8130, 6582, 6621, 5591, 5528, 7886, 6719, 6879, 7752, 7411, 7844, 8023, 7402, 10031, 10732, 9521, 9003, 11179, 4926, 0, 606, 0, 172, 0, 35, 0, 0, 0, 0, 0, 0, 0, 42, 0, 208, 0, 723, 0, 5933, 14090, 12046, 12678, 10625, 11458, 12280, 11967, 12215, 12495, 12428, 12805, 11910, 12014, 4610, 0, 265, 231, 0, 3884, 7180, 5598, 5525, 6440, 8057, 7469, 9286, 7943, 7233, 4772, 3984, 7659, 6953, 9917, 11242, 5205, 5562, 2460, 0, 163, 120, 0, 1016, 0, 8291, 17353, 14299, 13502, 10263, 8173, 5009, 5943, 5937, 6011, 5894, 5668, 6299, 7843, 7033, 9387, 12410, 12776, 13457, 13356, 13688, 12416, 11470, 8774, 10723, 5202, 0, 671, 0, 190, 0, 37, 0, 0, 0, 0, 0, 0, 56, 0, 277, 0, 962, 0, 7809, 17879, 14361, 16010, 15372, 15929, 16688, 16390, 16244, 15538, 15672, 14469, 14683, 11456, 9809, 9864, 11379, 12471, 8435, 10883, 11332, 8602, 6850, 4208, 807, 0, 48, 0, 12, 0, 43, 0, 200, 0, 701, 0, 5577, 12229, 9829, 10951, 10387, 10623, 10614, 10375, 11671, 14026, 9502, 5520, 6096, 6310, 6543, 6465, 6359, 6454, 5968, 4765, 9344, 12387, 12072, 13227, 13463, 13105, 13574, 12240, 9994, 6689, 1159, 0, 54, 0, 0, 20, 0, 173, 0, 614, 0, 5393, 14291, 12360, 12478, 13443, 13893, 13800, 13815, 13836, 13787, 13872, 13584, 13711, 15344, 13049, 10644, 11489, 11312, 11948, 9729, 7426, 7312, 6794, 6308, 6490, 2592, 0, 270, 0, 67, 0, 0, 195, 0, 740, 0, 4505, 3371, 2042, 9354, 4872, 745, 292, 0, 4169, 10219, 9676, 10769, 9499, 9173, 9255, 9142, 9328, 9008, 9615, 7612, 5348, 5847, 5561, 5670, 5337, 7396, 10494, 11632, 12321, 12327, 11960, 10486, 9461, 6914, 5898, 2560, 0, 322, 0, 89, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24827, 23303, 21950, 22786, 20071, 16554, 16800, 17476, 19474, 20910, 20768, 20371, 19778, 19996, 19855, 19988, 19810, 20125, 19125, 18487, 20552, 21755, 22457, 22488, 21724, 22007, 21899, 21103, 19447, 18111, 17828, 17104, 16129, 15885, 13925, 13028, 12748, 14914, 14828, 14631, 17414, 18153, 17668, 16519, 17123, 16591, 16910, 17477, 18190, 19466, 19424, 18263, 18827, 18889, 18738, 17942, 17017, 17345, 17121, 17344, 17038, 17592, 15717, 13137, 13350, 13288, 14711, 15532, 15241, 15922, 17759, 17513, 17027, 16313, 14782, 16010, 17884, 19209, 19166, 18752, 19238, 18287, 17753, 18779, 17398, 16140, 15374, 15049, 15084, 14534, 14207, 13428, 13692, 13844, 14660, 15865, 15827, 17142, 17267, 17997, 19125, 18749, 18949, 18825, 18922, 18811, 19007, 18572, 18444, 18820, 18758, 17606, 16181, 15532, 14839, 14921, 14745, 13761, 14331, 13996, 13650, 15786, 15597, 14792, 15538, 16410, 17164, 17854, 17662, 17186, 17149, 16269, 15603, 17068, 18357, 19056, 18867, 18346, 18646, 18059, 16174, 14646, 15182, 14877, 14308, 14529, 14344, 14568, 14233, 14854, 12775, 11004, 15370, 16194, 15996, 16733, 15586, 15462, 15382, 15220, 15682, 17931, 18526, 16855, 16536, 17467, 17580, 16827, 15608, 14875, 15149, 15197, 15142, 14573, 13679, 13817, 13585, 16570, 13020, 11703, 15809, 16023, 17942, 17006, 15872, 15009, 15649, 16021, 15633, 15766, 15730, 15687, 15825, 15520, 16522, 17239, 16186, 16092, 15926, 15980, 15647, 15429, 15728, 15524, 15411, 16644, 17510, 16475, 16691, 17746, 17492, 17348, 17271, 16667, 16801, 17214, 17979, 17314, 17281, 17412, 16858, 18022, 17753, 17189, 16884, 16971, 16815, 16577, 15935, 16460, 13154, 10154, 11166, 10617, 11022, 10603, 11195, 10116, 13574, 17003, 16029, 16676, 16931, 17873, 18292, 16908, 16128, 17049, 17442, 17379, 16897, 16693, 16863, 16609, 16562, 15597, 15953, 14110, 10783, 14439, 16741, 14763, 14519, 16059, 16006, 16236, 17788, 14913, 11276, 14571, 16497, 15780, 16010, 15917, 15122, 15226, 16134, 15860, 15930, 16023, 15717, 16420, 14142, 11948, 9747, 10037, 7910, 8384, 10295, 8443, 11440, 14620, 14366, 11060, 9647, 10079, 9848, 12391, 13321, 14063, 13087, 9878, 11550, 11823, 12439, 12216, 12425, 12403, 12889, 9611, 7884, 3186, 501, 8794, 5963, 6825, 9966, 7206, 10090, 11483, 11706, 11689, 11646, 11728, 11595, 11840, 11066, 10473, 11321, 11925, 12732, 12832, 12588, 12793, 12936, 12579, 9048, 5663, 5956, 4887, 6947, 6082, 3270, 4690, 5598, 4459, 6837, 8356, 6945, 8410, 8428, 9013, 8378, 9507, 10226, 9651, 10852, 11167, 11763, 12359, 12165, 11536, 12155, 11176, 9988, 10191, 10362, 9793, 11068, 6634, 1469, 2631, 0, 4397, 8443, 6219, 8214, 8255, 8533, 8033, 8797, 9642, 10100, 10470, 10673, 11268, 11390, 11518, 11321, 12483, 9601, 6598, 6575, 5978, 5504, 4422, 2128, 3414, 6290, 2386, 0, 2135, 3727, 4206, 6798, 7833, 7991, 9176, 10217, 9936, 10027, 10059, 9876, 10558, 11175, 11266, 10686, 8319, 6894, 6437, 5584, 5322, 3894, 4323, 6037, 6804, 2491, 58, 3134, 2978, 4151, 5035, 7151, 9500, 9024, 9962, 10352, 10040, 10397, 10341, 10341, 10404, 10634, 10406, 9529, 7279, 6453, 6682, 4878, 4217, 5452, 6377, 6647, 6551, 6636, 6539, 6697, 6084, 6269, 12636, 11962, 7771, 9714, 9645, 9700, 10704, 10949, 11130, 11117, 12570, 14430, 12682, 11310, 9426, 6969, 8344, 7955, 5929, 8512, 11145, 11638, 12830, 9050, 6437, 8008, 7705, 12367, 17315, 13801, 10400, 10538, 10193, 10652, 11114, 11546, 11758, 11733, 11664, 11867, 11441, 12302, 9900, 9526, 8517, 9647, 12835, 11665, 12375, 11715, 10319, 8431, 11811, 13302, 12969, 14470, 14157, 16623, 12793, 12638, 16974, 16295, 17045, 17155, 17427, 16993, 17986, 17635, 18901, 14693, 13401, 14770, 12255, 13531, 13139, 13854, 14355, 13797, 13457, 14363, 14795, 14664, 14776, 14625, 14873, 14397, 15949, 17580, 17203, 17482, 17761, 17670, 17172, 16817, 17327, 15629, 12998, 13460, 12791, 12873, 14604, 14022, 14842, 15320, 15041, 15680, 16200, 18144, 18809, 19861, 20653, 20053, 19106, 17950, 18014, 18050, 17567, 17819, 18205, 17803, 17581, 16678, 17546, 15124, 12454, 13238, 12924, 12946, 13207, 12510, 14890, 16942, 16187, 17452, 18525, 20475, 20669, 21861, 23046, 20743, 18435, 18242, 18625, 18320, 18427, 18462, 18227, 17624, 17648, 17062, 17353, 14548, 14667, 16540, 15683, 16641, 16974, 17680, 18527, 17415, 16881, 17541, 19798, 21595, 22813, 23696, 24534, 23016, 20474, 21337, 20839, 21220, 20803, 21471, 19389, 17086, 17423, 17280, 17093, 16928, 16849, 16643, 17718, 18656, 18534, 19413, 18627, 17502, 17742, 19650, 22648, 23893, 24843, 24916, 24590, 22090, 20280, 19545, 18644, 18508, 18704, 18809, 18151, 18085, 17696, 17771, 17198, 17263, 17959, 17860, 18175, 17714, 17531, 17509, 17637, 17357, 17904, 16790, 20479, 24503, 24378, 24587, 23577, 22278, 19938, 19175, 18926, 19180, 18880, 18260, 18440, 18004, 18202, 17612, 17340, 17669, 16886, 18174, 18950, 18117, 20330, 22900, 22404, 22436, 22918, 22894, 24443, 24045, 26825, 27457, 24345, 23626, 21789, 20434, 19142, 19289, 19376, 19379, 19341, 19428, 19257, 19617, 18366, 17069, 18375, 19608, 18228, 20173, 22260, 22409, 22910, 21841, 22929, 23644, 24278, 24919, 24719, 23349, 23038, 22568, 20837, 19486, 19419, 19712, 19330, 19654, 18709, 18306, 17537, 18007, 17913, 17260, 17903, 18104, 17783, 19337, 21521, 21800, 21047, 19612, 19697, 19577, 19686, 19547, 19769, 19350, 20634, 21165, 19399, 19670, 19704, 19600, 19726, 19118, 18479, 17702, 17938, 18820, 18447, 18259, 18499, 18520, 18582, 21639, 23615, 22550, 22238, 22914, 24269, 24755, 25429, 24643, 23740, 23593, 23522, 21675, 19453, 19386, 19457, 19869, 19504, 19435, 19773, 19235, 18942, 19009, 18986, 18980, 19023, 18888, 19635, 22379, 23567, 20222, 20910, 24485, 24989, 25582, 25528, 24606, 24014, 24534, 22598, 20480, 20445, 19985, 20138, 20314, 20066, 20147, 19942, 19432, 19639, 18914, 20280, 22017, 19227, 19966, 23602, 23832, 23524, 23317, 22470, 24124, 25479, 25833, 25897, 24635, 24365, 24444, 24317, 24550, 24126, 24962, 22192, 19222, 20022, 19690, 19733, 19586, 19573, 23109, 25458, 22408, 22667, 24978, 25280, 25021, 24659, 24339, 25284, 25096, 27837, 31847, 27329, 24092, 24183, 24023, 23099, 20579, 20129, 20568, 21501, 22379, 21341, 20269, 19426, 20745, 24142, 25689, 26055, 26294, 26526, 26480, 26459, 26547, 26369, 26704, 25874, 27474, 31306, 27604, 24390, 24367, 24171, 22117, 19854, 20281, 19907, 19839, 19958, 19911, 19695, 18999, 19510, 19382, 18701, 18633, 18516, 19149, 20946, 23617, 25632, 20049, 14693, 20981, 24792, 24513, 25090, 24236, 23936, 22501, 20499, 20050, 20006, 19768, 19545, 19610, 19580, 19595, 19587, 19598, 19552, 19241, 18624, 19089, 19559, 20370, 20814, 20221, 17408, 15032, 18503, 20929, 22213, 23487, 21605, 20467, 19909, 19494, 19773, 19454, 19228, 19555, 19132, 18893, 18928, 18641, 19097, 19252, 19557, 19452, 18135, 18300, 19125, 21738, 22734, 22983, 22385, 21535, 22534, 22117, 22361, 22181, 22366, 22074, 23026, 23913, 22071, 21859, 23328, 23669, 23257, 21374, 18858, 19278, 19475, 21967, 23877, 23584, 24448, 24066, 24719, 25345, 24815, 25084, 24319, 26742, 29924, 29007, 29994, 25845, 22544, 23261, 23849, 22853, 20958, 20823, 22158, 22873, 21023, 19182, 18002, 18148, 18098, 18069, 18201, 17918, 18447, 17392, 20949, 24996, 23167, 23673, 23023, 26825, 29637, 28928, 24533, 20936, 22738, 23083, 21612, 19343, 18532, 19661, 19326, 17602, 17961, 17696, 17826, 17698, 17333, 17624, 17666, 17670, 17897, 21190, 22599, 22498, 21166, 19308, 21406, 22619, 21759, 17562, 16025, 16996, 16931, 17013, 16980, 16967, 17029, 16888, 17331, 17563, 17434, 17697, 17926, 17817, 17229, 17121, 16715, 18702, 21546, 22063, 21399, 21715, 20350, 24263, 28108, 26433, 22960, 18727, 20421, 23169, 22991, 21050, 21796, 22737, 22395, 20909, 17732, 16648, 16945, 16414, 16237, 15959, 17581, 20243, 18955, 20546, 22597, 22073, 22140, 22461, 21555, 24680, 26869, 24259, 23947, 24418, 25476, 24521, 24360, 24982, 26431, 23929, 19826, 17183, 15730, 15623, 15452, 15397, 16692, 18690, 20923, 21835, 24304, 27950, 27941, 28385, 28043, 28227, 28976, 28720, 27647, 25687, 25126, 25696, 26375, 26261, 26689, 27291, 27152, 26689, 26044, 26115, 26335, 25746, 26990, 23505, 23793, 24912, 25250, 29163, 28727, 29931, 29741, 29221, 29529, 29811, 29946, 29309, 27901, 27387, 27662, 28351, 28098, 27919, 28656, 28386, 29614, 24436, 20148, 21068, 20011, 19685, 20412, 21642, 24067, 26700, 27541, 29830, 30234, 30400, 30631, 30389, 30530, 30796, 31050, 30934, 31054, 30886, 31180, 30217, 29083, 30646, 30151, 31673, 26606, 25234, 24882, 23584, 27685, 27120, 28938, 29383, 29507, 29909, 30394, 30803, 31030, 30737, 30945, 31046, 30907, 31280, 31082, 30718, 30545, 30680, 30936, 30525, 30818, 30831, 31431, 30577, 25618, 23762, 23249, 23274, 22954, 25565, 28172, 27415, 27715, 27697, 27421, 28540, 29289, 29556, 30693, 31116, 31764, 31850, 31239, 31041, 31519, 31586, 31512, 31432, 32021, 31986, 32023, 27614, 24881, 24625, 26050, 29213, 29185, 30939, 31359, 30585, 30627, 30197, 29774, 29864, 30005, 29775, 30790, 31996, 31599, 31594, 31884, 31727, 31609, 31644, 31689, 31555, 31823, 31320, 32343, 28785, 24415, 27153, 29545, 30404, 30854, 30444, 30369, 31092, 31164, 30679, 30775, 31211, 30958, 30969, 31496, 31928, 31598, 31175, 31987, 32559, 32465, 32757, 31076, 30084, 30792, 31434, 30637, 29171, 28432, 28696, 30293, 31410, 32059, 31820, 31090, 30875, 30871, 30689, 31087, 30261, 31781, 29043, 34431, 16233, 0, 4445, 0, 17111, 35683, 26620, 27639, 28032, 30647, 29491, 27740, 26493, 26408, 27611, 30635, 31939, 31178, 29315, 29867, 29652, 29003, 29351, 29827, 28935, 30592, 29688, 35160, 18370, 0, 18131, 34765, 30585, 30698, 27020, 27639, 27141, 27423, 27325, 27341, 27345, 27325, 27360, 27298, 27599, 28415, 27552, 27562, 27036, 28992, 29157, 26337, 27206, 26419, 29263, 32019, 31766, 32253, 29820, 27920, 28436, 27450, 25834, 25101, 25715, 26420, 26237, 26146, 25779, 25869, 26198, 27280, 27924, 27445, 27351, 27108, 26811, 27801, 27257, 25963, 26075, 26262, 26500, 26413, 26471, 26407, 26504, 26355, 26398, 23337, 20508, 22219, 24124, 25138, 23782, 22983, 24673, 25549, 26448, 27348, 27265, 27296, 26384, 26429, 27255, 27149, 26483, 26608, 26797, 27500, 28324, 28251, 28753, 27758, 27364, 27214, 26853, 21151, 17309, 18027, 18295, 20655, 20893, 21673, 21766, 23432, 25104, 24570, 24864, 24659, 24852, 24569, 25449, 26468, 25817, 25610, 27018, 28145, 28020, 27835, 27285, 27125, 26234, 24478, 22669, 18654, 18324, 18751, 19930, 19568, 18064, 17750, 19933, 22847, 24589, 24924, 23090, 24048, 23357, 24647, 25336, 24932, 23879, 24609, 26367, 26326, 26988, 26812, 25879, 24885, 24547, 24702, 24487, 24848, 24206, 25468, 21344, 17155, 18102, 17371, 21763, 25346, 22727, 23152, 24405, 23627, 24967, 24497, 24611, 23449, 24166, 24743, 25163, 26087, 25211, 24759, 23473, 23779, 20698, 18200, 17226, 17106, 18335, 18484, 16242, 16934, 14934, 15767, 21102, 21040, 22929, 22737, 22154, 23626, 24312, 24149, 24243, 24154, 24271, 24068, 24652, 24808, 24267, 23293, 23515, 20828, 18506, 17863, 17808, 18819, 18705, 16798, 15493, 17209, 17133, 19760, 22135, 22748, 23389, 22771, 22483, 24381, 24358, 23552, 23616, 24152, 23963, 23308, 24362, 24299, 23978, 23136, 21977, 19440, 18322, 17576, 17633, 18487, 18024, 18206, 18158, 18104, 18273, 17884, 19490, 22395, 20822, 21774, 25095, 23043, 23001, 23426, 23051, 23526, 23680, 24462, 24158, 23090, 22170, 22735, 20110, 18091, 18859, 18071, 18186, 18856, 19203, 20082, 18806, 18907, 20476, 21502, 20430, 21055, 22833, 22860, 23352, 22815, 23343, 23239, 22957, 22711, 22430, 22574, 22406, 22671, 22204, 23121, 20212, 17755, 18547, 18257, 18461, 18541, 19607, 17083, 17891, 20323, 21007, 20876, 22086, 22410, 22817, 24255, 23612, 23526, 22754, 23120, 22708, 23187, 24257, 23706, 22752, 23266, 22201, 19259, 18297, 18219, 17103, 17127, 17183, 19308, 19908, 18547, 19506, 19892, 20249, 20106, 20219, 20076, 20311, 19859, 21273, 22515, 22633, 23245, 22632, 23815, 23911, 22521, 22401, 20073, 18120, 18054, 18014, 17814, 17971, 18165, 18537, 16564, 15180, 17892, 20401, 18504, 18729, 22832, 22055, 23042, 22697, 20864, 21114, 21579, 22934, 23016, 23556, 23841, 22363, 21534, 19708, 18540, 18904, 18779, 18754, 18935, 18529, 19389, 16435, 13695, 18224, 20824, 18701, 19047, 21747, 22007, 22646, 21512, 21715, 23226, 23368, 24220, 23546, 23473, 23762, 22753, 22957, 20355, 18551, 18405, 18033, 18316, 17892, 18295, 19000, 18490, 15533, 16486, 19454, 19697, 17963, 19291, 21022, 22233, 21792, 20349, 21132, 20779, 20960, 20878, 20896, 20923, 20903, 21317, 19922, 18181, 17921, 18008, 18019, 17998, 18272, 18762, 16893, 14563, 16807, 18937, 17422, 16225, 19268, 21363, 21424, 20372, 19749, 20813, 21611, 22818, 23386, 23281, 23690, 22051, 20692, 19504, 18409, 18730, 17939, 18206, 18433, 17192, 15322, 13117, 12240, 12388, 12454, 12170, 12783, 11498, 15723, 19775, 18987, 19126, 20895, 22353, 22079, 23464, 22999, 23698, 22383, 21241, 19563, 17989, 18364, 17897, 18097, 17802, 15213, 13288, 12418, 13422, 15746, 17265, 17545, 17782, 17214, 18398, 19881, 19464, 19375, 20848, 23091, 22985, 23480, 23249, 23586, 22805, 21953, 22143, 22168, 21942, 22504, 20374, 17394, 18274, 15260, 13870, 17311, 17943, 19108, 19138, 18143, 17238, 20752, 23949, 22374, 23700, 24640, 24624, 24346, 24014, 23609, 23281, 23067, 23145, 23801, 22204, 19590, 18430, 18265, 18690, 18674, 19249, 19434, 19172, 18678, 19310, 20710, 21874, 21192, 21873, 23283, 22834, 23039, 22968, 22916, 23401, 24789, 25139, 24943, 24554, 24020, 24410, 23126, 22304, 20421, 19779, 20679, 21223, 21568, 20706, 20731, 19920, 22565, 25267, 24609, 24300, 24851, 25946, 26147, 26082, 26435, 26154, 26036, 25472, 25724, 26009, 25443, 24488, 24474, 24559, 23260, 20319, 20752, 20653, 18766, 19555, 18946, 19637, 18513, 22076, 26322, 25213, 25718, 25993, 26885, 27463, 27484, 27677, 27026, 26653, 26006, 26174, 26651, 25916, 25138, 25057, 24872, 24043, 23790, 23974, 23413, 23839, 24710, 24651, 23727, 23418, 25067, 25722, 25569, 25742, 26195, 26377, 27095, 27118, 27225, 27558, 27097, 26315, 25824, 25924, 25949, 25801, 26149, 25024, 23987, 23193, 22049, 23018, 23247, 24997, 25008, 23339, 24567, 25334, 25354, 25578, 25991, 26430, 26305, 26734, 27097, 27317, 27295, 26701, 26225, 26137, 26711, 26157, 25947, 25367, 25368, 24770, 23278, 20231, 18775, 19229, 20506, 22145, 21923, 21223, 22478, 24209, 23629, 23981, 23681, 24043, 23426, 25448, 28000, 27322, 26942, 26282, 26321, 27415, 26961, 25716, 25716, 24885, 25597, 14476, 2420, 0, 2925, 7566, 8640, 7839, 6278, 7122, 2919, 0, 145, 0, 25, 19, 0, 222, 0, 771, 0, 6494, 15692, 12175, 17745, 21100, 19680, 20392, 20392, 22325, 31593, 28643, 37154, 11462, 12254, 38560, 28409, 32570, 29652, 29482, 30316, 32696, 32029, 31416, 30564, 28882, 27659, 27538, 27313, 27168, 27368, 27338, 28684, 28413, 32110, 27506, 36466, 14197, 8308, 30218, 23915, 27328, 25665, 26196, 26641, 23720, 19127, 18894, 22034, 24441, 26333, 13012, 1580, 4898, 5081, 6648, 6750, 7238, 6036, 6012, 6187, 5095, 4729, 4679, 5481, 4469, 3951, 3050, 1209, 1099, 1134, 809, 1524, 1138, 345, 493, 0, 869, 1728, 440, 0, 30, 0, 10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 60, 0, 210, 0, 1957, 5729, 5045, 9883, 16043, 20195, 22489, 21688, 22315, 21565, 22725, 20555, 27324, 32319, 28490, 30073, 29136, 25827, 24024, 22032, 22276, 11781, 3339, 11149, 19106, 14785, 10923, 7345, 1159, 1530, 233, 1582, 1272, 1595, 1007, 519, 1399, 2767, 3362, 3279, 3918, 4383, 4287, 4744, 4865, 4405, 4250, 3967, 3888, 3029, 2380, 2563, 2486, 2501, 2544, 2396, 2905, 3223, 3475, 2849, 4143, 1766, 9298, 18151, 23108, 11139, 0, 1823, 0, 2298, 4262, 5673, 10226, 4165, 0, 485, 0, 147, 0, 32, 0, 0, 0, 0, 0, 15, 0, 76, 0, 266, 0, 2342, 6481, 6827, 7356, 7002, 7434, 6748, 7956, 5566, 13469, 22020, 20282, 21319, 20336, 20625, 20359, 20074, 21325, 22512, 21183, 20033, 19334, 18340, 18172, 17867, 17180, 17079, 17499, 17614, 18298, 18932, 20933, 19250, 16906, 11811, 8660, 10461, 9696, 7935, 7189, 7653, 8029, 7397, 1846, 25, 5143, 11253, 12787, 12629, 12429, 13007, 11837, 14238, 6307, 0, 780, 0, 220, 0, 22, 192, 1481, 2239, 1568, 405, 0, 364, 2371, 2957, 1309, 565, 112, 0, 10, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 261, 2076, 2985, 2387, 2221, 0, 7152, 16726, 15195, 16513, 16069, 16050, 15787, 14898, 14910, 16278, 5446, 0, 2970, 3140, 4633, 5102, 5224, 5260, 5122, 5401, 4895, 5899, 2610, 0, 324, 0, 92, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 31, 0, 100, 0, 937, 2615, 1768, 3437, 4896, 4519, 4614, 4732, 4353, 5208, 2312, 0, 286, 0, 82, 0, 27, 0, 55, 0, 258, 0, 1598, 661, 734, 0, 8917, 20743, 20125, 23821, 23065, 24738, 26154, 27185, 28283, 29741, 30523, 31892, 31776, 31309, 31981, 30335, 28804, 28416, 27885, 27292, 25332, 22013, 20339, 20837, 20501, 20850, 20368, 21224, 18425, 15329, 17639, 17358, 21210, 20655, 17070, 18594, 17951, 16012, 13861, 14021, 16189, 18016, 19676, 20122, 23352, 26653, 21639, 23850, 9490, 0, 3682, 1353, 2630, 1637, 2495, 1528, 463, 684, 516, 221, 0, 0, 92, 0, 896, 2181, 1926, 2096, 1962, 2108, 1894, 2291, 1013, 0, 125, 0, 36, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 79, 0, 284, 0, 3847, 12321, 17497, 18691, 18993, 19304, 20021, 20116, 19060, 19106, 15165, 20847, 19844, 4360, 0, 1865, 3924, 4853, 5370, 5579, 6221, 4473, 3543, 1365, 0, 160, 0, 24, 15, 0, 266, 266, 0, 51, 0, 13, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 35, 0, 103, 0, 1089, 3358, 1629, 6004, 10322, 9379, 9274, 9762, 14890, 17807, 20562, 15978, 3130, 0, 188, 0, 61, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 93, 0, 458, 0, 1596, 0, 13195, 31663, 27884, 30856, 30795, 31810, 31834, 31989, 31762, 31887, 30204, 28494, 26426, 24549, 24301, 23658, 23802, 23970, 23932, 21425, 19260, 18702, 18642, 18142, 18912, 21306, 21038, 20941, 21333, 22113, 21593, 22521, 19384, 17258, 19322, 18741, 18853, 18118, 18117, 17914, 18336, 17535, 19016, 16096, 25485, 32040, 19062, 15604, 13517, 15914, 8336, 13, 1153, 0, 399, 0, 76, 0, 8, 0, 12, 0, 52, 0, 183, 0, 1607, 4486, 4369, 3972, 3103, 4021, 1738, 0, 214, 0, 61, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 4, 0, 16, 0, 144, 287, 138, 748, 1922, 2082, 1442, 1751, 0, 7004, 18375, 19209, 23959, 23854, 26913, 30152, 29048, 29767, 29071, 30112, 26717, 18395, 4432, 1601, 6018, 13486, 12716, 5813, 7022, 1407, 0, 152, 0, 1175, 2207, 2108, 2709, 2943, 3861, 4174, 3989, 4313, 4399, 4100, 3718, 3799, 3487, 3373, 3378, 3285, 2436, 2717, 3334, 2616, 2846, 2918, 2840, 2474, 2916, 3529, 3332, 3414, 3406, 3388, 2983, 895, 7415, 15036, 14340, 20465, 20615, 5320, 0, 443, 0, 135, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 14, 0, 57, 0, 1365, 8805, 17454, 26433, 31537, 31205, 32117, 32674, 32617, 32599, 32531, 32642, 32421, 32832, 32071, 33599, 28587, 23536, 24825, 24813, 24022, 22063, 21186, 19272, 18643, 18552, 18418, 17065, 16663, 11417, 5260, 5506, 5862, 7392, 10112, 10297, 8979, 9004, 9735, 9744, 10173, 9181, 8302, 6846, 6067, 4183, 1432, 0, 4305, 5378, 1765, 3988, 3732, 1925, 0, 308, 0, 130, 32, 88, 27, 0, 3, 0, 8, 0, 30, 43, 1240, 2681, 4701, 5476, 3655, 4085, 1737, 0, 214, 0, 62, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 45, 0, 162, 0, 1122, 1476, 380, 194, 168, 0, 1018, 0, 8714, 21222, 20499, 22482, 26498, 30915, 31044, 30654, 31987, 28271, 23229, 20028, 5415, 0, 1623, 3158, 12203, 12131, 8920, 7985, 912, 17, 0, 5, 5, 0, 4, 0, 0, 10, 0, 41, 0, 304, 598, 1148, 1774, 2721, 3647, 3872, 3923, 1201, 0, 121, 0, 35, 0, 1, 7, 0, 42, 0, 390, 1269, 1593, 1834, 1736, 2342, 1907, 4006, 8196, 2898, 0, 742, 0, 164, 0, 41, 0, 3, 0, 0, 0, 0, 0, 4, 0, 0, 23, 0, 331, 1042, 2734, 0, 12011, 28882, 21510, 21134, 21317, 22922, 24615, 25016, 26695, 26763, 26303, 26341, 26302, 26160, 26485, 26042, 27062, 28192, 27100, 26568, 21934, 18580, 17780, 16690, 16721, 15408, 14913, 15121, 14836, 15319, 14467, 16139, 10681, 5516, 8732, 7910, 7929, 8724, 9810, 9531, 9371, 9526, 7566, 2113, 19733, 31309, 22662, 19571, 17335, 18761, 16518, 14958, 15034, 5561, 0, 854, 0, 198, 0, 51, 0, 24, 0, 63, 0, 886, 3636, 2478, 1659, 2762, 2538, 2718, 2566, 2743, 2472, 2984, 1320, 0, 163, 0, 46, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 9, 0, 31, 0, 256, 575, 483, 518, 518, 483, 575, 256, 0, 31, 0, 3, 6, 0, 35, 0, 252, 282, 0, 94, 0, 898, 4176, 3671, 553, 0, 10, 0, 4, 0, 0, 2, 0, 28, 0, 100, 0, 866, 2237, 2197, 2532, 3106, 3446, 3566, 3837, 3804, 3850, 3788, 3885, 3717, 4056, 2797, 1168, 4002, 6591, 6040, 5532, 7782, 7230, 9757, 11451, 10191, 13035, 13872, 9570, 6408, 7011, 4697, 4607, 2249, 705, 1575, 143, 26, 0, 3, 0, 0, 1, 0, 56, 0, 297, 0, 1063, 0, 8698, 21504, 24852, 29497, 28136, 28251, 29284, 26682, 32239, 14743, 993, 169, 14286, 32428, 26204, 28683, 26776, 27276, 26654, 26499, 26291, 26398, 25976, 25716, 25347, 25146, 25370, 25398, 26151, 25376, 26359, 23119, 19166, 19800, 19938, 19316, 18578, 19052, 18915, 19543, 20100, 20066, 19618, 21096, 20846, 21241, 22555, 21917, 22432, 21760, 22848, 20934, 24707, 12257, 0, 3228, 1342, 2549, 1004, 170, 536, 0, 1129, 2035, 175, 3050, 4895, 3320, 1484, 571, 2317, 2434, 3993, 4533, 4784, 3511, 328, 21, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 22, 0, 63, 0, 779, 3246, 3179, 5058, 5672, 11622, 16810, 15168, 15022, 14483, 13498, 13484, 3006, 5049, 19762, 21699, 26275, 29318, 30637, 29894, 28776, 29274, 28784, 29474, 28303, 30573, 23323, 16761, 18506, 18096, 18017, 15032, 16094, 15459, 17656, 11036, 5592, 7130, 7245, 4846, 1236, 2689, 2268, 2343, 2013, 2693, 2339, 3764, 753, 8480, 17301, 17301, 18935, 18567, 20391, 20115, 20990, 22571, 26746, 28270, 26981, 28335, 28823, 29233, 29807, 29441, 29950, 29090, 30566, 27931, 33830, 18536, 0, 18678, 33652, 27199, 26685, 27533, 14108, 0, 780, 0, 220, 0, 32, 0, 0, 42, 0, 117, 0, 1338, 4463, 2589, 9530, 16306, 20159, 25518, 29156, 32114, 31116, 31210, 30531, 29944, 29742, 29668, 29409, 29263, 29098, 29030, 29277, 28765, 29852, 26091, 21517, 21790, 21525, 17936, 17986, 10731, 4170, 7933, 8008, 8999, 9255, 9685, 9784, 10449, 10508, 10477, 10713, 9571, 8755, 9197, 9187, 9146, 8807, 8113, 7591, 6808, 6973, 6244, 3682, 1126, 1396, 1513, 0, 668, 1089, 420, 47, 0, 9, 0, 28, 0, 100, 0, 1104, 4277, 5578, 3355, 1313, 986, 155, 0, 3, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 58, 0, 266, 0, 2035, 3875, 5498, 2632, 13344, 26776, 25892, 28569, 28298, 27999, 29193, 25097, 21171, 22638, 26916, 29437, 29205, 26063, 26496, 11051, 0, 3271, 5819, 12136, 15533, 17774, 16242, 17204, 19171, 9821, 2019, 4354, 3243, 3761, 3637, 3410, 4117, 1714, 0, 0, 1995, 5137, 3537, 2735, 2541, 2477, 2788, 2588, 2919, 3548, 3051, 964, 513, 895, 737, 969, 173, 72, 0, 723, 988, 668, 377, 1959, 3558, 3929, 6491, 3728, 1126, 1316, 1361, 728, 0, 96, 0, 23, 0, 4, 0, 0, 0, 0, 3, 0, 50, 0, 228, 0, 1850, 5602, 16353, 23943, 27347, 28480, 36249, 16609, 0, 1339, 1719, 0, 15635, 37745, 28970, 36844, 18079, 0, 17744, 33334, 28242, 29498, 26746, 25090, 23679, 22940, 23057, 23285, 22878, 22050, 21673, 21931, 21917, 21756, 22152, 21373, 22937, 17928, 13722, 15518, 13812, 14643, 13514, 14810, 19277, 21035, 21522, 19224, 21807, 10272, 0, 2949, 190, 14, 327, 788, 544, 556, 581, 263, 0, 16, 8, 0, 88, 0, 1020, 3869, 5401, 6546, 6966, 4503, 3127, 1313, 0, 168, 0, 46, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 29, 0, 105, 0, 694, 694, 0, 105, 0, 29, 0, 2, 2, 0, 19, 0, 70, 0, 743, 2740, 4069, 4904, 5101, 2966, 2254, 1191, 0, 165, 0, 45, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 54, 0, 194, 0, 1273, 1273, 0, 194, 0, 54, 0, 10, 0, 0, 0, 0, 9, 0, 43, 0, 150, 0, 1217, 2720, 1694, 551, 0, 63, 0, 15, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 103, 0, 252, 0, 3600, 17736, 22107, 32504, 15737, 0, 2424, 101, 473, 1912, 0, 12472, 27248, 22810, 25556, 24510, 24979, 25042, 25059, 24749, 24619, 23618, 23617, 23925, 23555, 22951, 22080, 21681, 20947, 20579, 18717, 17273, 17656, 16591, 14548, 13167, 14036, 14633, 14402, 14348, 13925, 9286, 8254, 6380, 9273, 2677, 7468, 8754, 0, 1778, 0, 860, 387, 556, 578, 271, 47, 430, 171, 0, 4, 20, 0, 61, 63, 1406, 2877, 723, 6107, 0, 21350, 20420, 0, 3098, 0, 875, 0, 168, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 55, 0, 202, 0, 1472, 2964, 3732, 4091, 780, 0, 35, 0, 0, 1732, 14544, 23468, 24931, 27062, 26445, 29073, 26695, 25117, 9377, 0, 1241, 852, 3029, 2672, 2891, 2894, 2634, 3301, 1985, 4234, 0, 12960, 11935, 0, 1798, 0, 507, 0, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 7, 0, 28, 0, 221, 703, 1171, 1971, 1663, 2587, 910, 7388, 12427, 11004, 10330, 14469, 19344, 18015, 18290, 18836, 17275, 20704, 9184, 0, 1139, 0, 0);

--  Datos (voy sustituyendo y ya, si no es inviable)
--    type t_reg_datos is array (0 to 32783) of integer range 0 to 30000;
    type t_reg_datos is array (0 to 30734) of integer range 0 to 30000;
    signal reg_datos_debug : t_reg_datos := (17166, 18722, 17136, 19328, 16272, 30682, 25392, 19056, 18718, 19600, 28924, 25336, 30720, 29354, 30166, 31610, 41556, 18268, 0, 10662, 23014, 25600, 26458, 26860, 27512, 26976, 26494, 26020, 28736, 24742, 24960, 24588, 20512, 20614, 20432, 26768, 29820, 30238, 30794, 30766, 28022, 26766, 27592, 27836, 27782, 27832, 27752, 27922, 27024, 23402, 20858, 21748, 25176, 25686, 26176, 27890, 29210, 30220, 29138, 30804, 28058, 24514, 23356, 22902, 20424, 16810, 9374, 11320, 20570, 16410, 16964, 12652, 0, 8194, 22212, 3974, 13850, 9938, 5560, 34044, 18020, 1996, 0, 5644, 20078, 17172, 13262, 14528, 13584, 14628, 13142, 15840, 7114, 0, 1546, 428, 0, 544, 0, 3816, 3296, 0, 0, 2572, 0, 18476, 21974, 20464, 27984, 0, 11898, 9018, 10686, 17864, 18054, 8342, 9228, 24354, 5704, 264, 970, 12992, 9768, 0, 15220, 20960, 21638, 23278, 27652, 27860, 26552, 27404, 26152, 28380, 24240, 32336, 9638, 8408, 10928, 686, 7042, 20064, 26814, 4570, 10814, 12110, 11536, 26152, 31052, 19482, 14126, 13928, 19376, 22004, 26876, 29814, 31054, 34062, 32506, 29940, 26598, 28698, 25864, 19364, 14890, 11806, 10506, 6660, 114, 3198, 4718, 0, 6746, 9468, 4638, 6346, 5586, 5766, 6108, 4990, 9350, 16158, 17828, 19206, 8304, 0, 10032, 22224, 22198, 24778, 21176, 18554, 3348, 6890, 24578, 16096, 14742, 14698, 12868, 13392, 10530, 16430, 17848, 9182, 14804, 17602, 11126, 0, 12102, 10082, 2888, 17568, 17126, 16716, 10012, 14258, 16584, 15042, 13576, 13868, 13932, 13540, 14398, 12560, 19354, 30922, 32954, 33514, 33322, 33268, 34874, 34986, 34920, 33760, 33272, 30552, 26686, 25614, 26384, 19446, 7714, 5780, 6592, 5994, 9846, 16552, 17776, 19762, 22286, 18290, 18372, 23914, 30388, 34542, 33950, 35382, 35218, 34616, 34734, 34430, 33354, 33300, 33692, 33658, 33522, 33854, 33232, 34494, 29728, 22726, 27876, 16900, 3710, 4424, 4348, 4522, 8754, 10304, 16692, 20644, 30518, 29280, 18118, 21800, 24398, 20804, 19886, 15072, 9110, 6040, 0, 1654, 0, 7650, 16150, 24838, 12958, 3610, 20516, 22354, 24372, 30912, 35082, 37306, 34808, 30654, 32524, 31906, 31754, 32716, 30608, 34950, 20858, 9964, 23124, 23434, 24332, 18144, 14018, 15036, 16420, 17966, 22678, 23168, 19812, 22624, 32658, 14580, 3056, 20162, 21830, 25550, 29600, 33116, 33644, 34424, 36744, 37322, 37376, 36116, 34232, 36446, 32980, 31954, 35916, 34752, 38054, 34980, 34980, 37450, 35404, 36246, 35894, 35892, 36234, 35446, 37070, 31618, 26406, 28398, 25490, 27872, 30224, 30588, 31832, 34702, 37246, 35840, 35926, 32574, 34978, 34376, 34464, 29976, 24310, 8874, 9036, 29194, 18044, 17416, 15258, 8388, 11428, 28268, 23460, 7838, 27976, 32574, 28330, 10028, 1148, 14780, 20444, 20012, 16434, 17718, 16950, 17572, 16904, 17938, 13880, 4848, 10860, 328, 9808, 6710, 8696, 23560, 0, 9688, 7086, 0, 1586, 20958, 26126, 12006, 15186, 22086, 11982, 0, 1504, 0, 524, 5642, 19918, 6546, 2998, 6602, 9014, 15208, 15498, 14868, 15588, 22668, 23314, 23766, 25432, 23884, 19268, 20532, 20484, 19394, 22030, 16630, 31216, 24794, 10544, 20830, 11668, 16954, 13182, 31704, 23266, 22766, 31160, 24804, 35322, 31824, 30072, 25514, 29162, 30742, 33156, 33864, 36512, 36858, 36478, 36448, 36364, 37094, 34724, 34180, 23958, 21760, 20900, 5256, 7114, 0, 7534, 8254, 5894, 10452, 3280, 5654, 5444, 3626, 8130, 0, 25206, 21434, 0, 1780, 4434, 18910, 17556, 19782, 17002, 18346, 4594, 5430, 12860, 5580, 13446, 16358, 17600, 14320, 21754, 17830, 16126, 12074, 11404, 14800, 4976, 1934, 2700, 15344, 13584, 0, 10182, 18626, 5074, 22568, 25186, 16182, 18768, 16534, 17948, 17096, 17806, 16924, 18356, 15552, 24954, 35964, 34392, 36296, 35718, 36434, 35636, 37196, 32736, 34470, 31582, 32938, 32174, 27362, 18572, 18048, 16346, 3570, 12446, 21476, 25554, 21702, 20982, 19276, 19924, 23028, 26776, 32058, 35010, 36286, 35970, 36738, 37086, 36568, 34768, 34072, 31978, 31952, 33962, 33472, 33318, 34138, 32354, 36068, 23584, 10054, 14098, 13922, 15768, 9356, 5660, 20088, 29218, 30760, 34806, 34636, 18716, 17010, 25488, 23560, 27658, 34048, 19070, 7716, 5494, 0, 1036, 910, 17864, 25510, 33392, 18756, 13798, 30138, 27904, 32986, 33012, 35632, 36598, 33498, 33400, 32596, 30576, 31246, 30938, 31028, 31134, 30754, 32126, 33892, 34914, 31276, 28600, 29984, 27148, 26052, 22902, 29112, 33560, 30244, 28424, 33270, 20400, 0, 8916, 22012, 26896, 31364, 31970, 32556, 31010, 33358, 33486, 32022, 32622, 30846, 32018, 32434, 35288, 38352, 37380, 39126, 37394, 35340, 34428, 31540, 31118, 31278, 30934, 31602, 30288, 34298, 36158, 31758, 32358, 28544, 28688, 31182, 31910, 34478, 35674, 35550, 35044, 34642, 33408, 33932, 34610, 29040, 37094, 16316, 19362, 14112, 3098, 23102, 22414, 9628, 2440, 27954, 34438, 37438, 34694, 28186, 27310, 21106, 14930, 16588, 13088, 26776, 30572, 19278, 22440, 20388, 21958, 20274, 22940, 15424, 12446, 13658, 10690, 1114, 6686, 6944, 2774, 23934, 11920, 14628, 11194, 0, 30144, 24112, 9482, 16764, 12874, 12294, 13268, 7772, 0, 11628, 4718, 9380, 10202, 2776, 10484, 0, 8798, 10544, 24546, 21340, 13136, 26192, 25596, 28396, 29264, 23466, 17824, 19746, 18466, 19674, 17892, 25328, 41126, 18866, 21460, 37406, 35618, 32460, 10064, 28876, 28042, 13142, 17464, 26166, 36082, 34516, 36666, 38676, 33204, 27830, 32192, 34246, 36164, 35860, 35478, 33224, 31594, 19530, 15750, 26126, 19622, 5428, 28036, 14984, 12096, 8486, 7184, 3984, 17234, 22882, 0, 4168, 0, 2696, 0, 15756, 40584, 21764, 15440, 14658, 9692, 25844, 35680, 32782, 35820, 23592, 3522, 0, 0, 2454, 13080, 16022, 11284, 16822, 10942, 0, 12790, 6322, 8082, 14348, 0, 11716, 9846, 0, 7910, 9146, 0, 4106, 0, 8486, 15540, 12536, 17780, 14706, 16030, 15576, 15392, 16230, 14278, 21282, 31514, 32616, 34160, 35094, 35274, 36012, 37094, 36602, 36882, 37114, 34336, 26906, 28006, 26294, 27606, 24634, 7032, 20930, 33176, 30940, 35334, 29858, 17942, 20682, 25448, 22216, 28828, 32604, 33842, 35576, 35752, 38188, 39192, 40028, 41040, 39076, 38284, 38296, 38330, 38250, 38378, 38200, 38540, 36432, 30238, 36122, 19430, 4076, 6922, 5792, 4192, 13762, 23536, 27898, 37856, 36904, 28610, 13210, 22604, 33962, 33902, 26428, 15332, 16332, 13370, 10808, 4278, 0, 4474, 23518, 28836, 36574, 14512, 4032, 26368, 24696, 32328, 29442, 29960, 32276, 23322, 19436, 20432, 19704, 20570, 19230, 21704, 14364, 9588, 11472, 22474, 34986, 29826, 28590, 29108, 19598, 9458, 12374, 12292, 10178, 20116, 28158, 23092, 3694, 6450, 22734, 27540, 32700, 33930, 34636, 34732, 36990, 37916, 38030, 38752, 35918, 32654, 36062, 37458, 37852, 36804, 40852, 35728, 33192, 38142, 35908, 36992, 36452, 36660, 36684, 36448, 37028, 35352, 32792, 31488, 28534, 29946, 32342, 33210, 34732, 35356, 36030, 35706, 35776, 34156, 34356, 32974, 34836, 30244, 34602, 5262, 18516, 22260, 3600, 30906, 11198, 7530, 18242, 14098, 27726, 25054, 13892, 16622, 15020, 9416, 10744, 14842, 25702, 38998, 35068, 37392, 35554, 37616, 34598, 40028, 23464, 10750, 13128, 0, 23160, 19736, 0, 3280, 25358, 8568, 17218, 22358, 0, 30870, 32902, 37406, 26742, 11134, 15582, 6784, 8734, 12192, 4034, 22596, 20948, 18214, 11102, 0, 8234, 12028, 19968, 16006, 13128, 25882, 26496, 29408, 30386, 29976, 28876, 29198, 29056, 29130, 29078, 29110, 29712, 34430, 32990, 35324, 38352, 42962, 24198, 24508, 39570, 31298, 37068, 34884, 34794, 36616, 37898, 38998, 33650, 30030, 29752, 31282, 34216, 34788, 33052, 32200, 26456, 23980, 27808, 16456, 5150, 32880, 20100, 5044, 8220, 0, 2478, 3342, 27144, 13570, 0, 1578, 0, 0, 916, 0, 8288, 14728, 15078, 8064, 1940, 28668, 26358, 14324, 20778, 8582, 0, 2706, 0, 14092, 24580, 9624, 2284, 980, 0, 11802, 8568, 4346, 9236, 0, 2442, 0, 1758, 0, 9336, 17694, 14926, 9576, 0, 9006, 4938, 4234, 15390, 13660, 16640, 15192, 16158, 15256, 16496, 14192, 21898, 31358, 30498, 32100, 34626, 35704, 33706, 31928, 33418, 29316, 29960, 27568, 18366, 25878, 21214, 13132, 14884, 13632, 16370, 24920, 34988, 37724, 32040, 32380, 27744, 28100, 34624, 33150, 34990, 35140, 36596, 39404, 40458, 39636, 40222, 40046, 38764, 37634, 36728, 37252, 36538, 37742, 35574, 39900, 25500, 9218, 11548, 13964, 14662, 13610, 20440, 20126, 27610, 32276, 33812, 3294, 18670, 27116, 11270, 37568, 22384, 14796, 10062, 6680, 4162, 0, 374, 2900, 22598, 28340, 34496, 14934, 2042, 23538, 19198, 26956, 30750, 32228, 27396, 27592, 20042, 21920, 36172, 31254, 33666, 32546, 32830, 33288, 30980, 28894, 29870, 29216, 29462, 29146, 26900, 27508, 19196, 8918, 15944, 23054, 26680, 20832, 1674, 7022, 22566, 26880, 31200, 32420, 34202, 33918, 35402, 35676, 35174, 34064, 30694, 28866, 31226, 32732, 34588, 37710, 39642, 39216, 38044, 37566, 33922, 32392, 32242, 32260, 32260, 32234, 32284, 32280, 30910, 21086, 18890, 25904, 27362, 30594, 33550, 34424, 33988, 32332, 32666, 29710, 26924, 29622, 31758, 28360, 18708, 10304, 15628, 15460, 9556, 18316, 6696, 2372, 14956, 10870, 22678, 34586, 35130, 25166, 11584, 13844, 16628, 15126, 28554, 37796, 38958, 29746, 19572, 22838, 21108, 22200, 21324, 22330, 19646, 16278, 17308, 3002, 2544, 0, 20804, 18748, 590, 15750, 0, 25154, 16570, 10412, 40788, 27476, 21696, 15066, 17600, 12346, 976, 5780, 19492, 18934, 18358, 20396, 18032, 24754, 31834, 24444, 2466, 9236, 20090, 19250, 22848, 25684, 24116, 27068, 36900, 33546, 35238, 34344, 34754, 34686, 33972, 26288, 6040, 5292, 17516, 14900, 28440, 29968, 29130, 35850, 32062, 33108, 32818, 35158, 36894, 32620, 25712, 26806, 31346, 29692, 31824, 23306, 27524, 25746, 8100, 14590, 9756, 18192, 6024, 8088, 11724, 0, 1236, 332, 0, 8846, 9180, 0, 1386, 0, 374, 0, 8, 80, 0, 350, 0, 3966, 15672, 17732, 18240, 17438, 18676, 7704, 0, 720, 2692, 18022, 4958, 6864, 12098, 0, 12396, 9730, 0, 1384, 0, 286, 92, 0, 1122, 0, 7666, 9542, 7104, 5598, 0, 306, 8280, 14670, 14702, 14686, 10272, 12086, 10802, 12142, 10026, 16970, 27398, 27780, 28906, 31264, 33750, 34788, 34684, 33140, 31786, 30438, 26748, 32674, 30576, 27758, 21312, 18270, 28066, 31538, 32584, 29102, 32676, 27024, 24462, 22014, 23278, 31276, 30610, 32178, 33320, 34872, 35182, 35634, 36220, 37744, 38756, 38672, 37100, 36804, 38134, 37352, 38334, 36696, 39754, 32136, 34500, 20318, 3036, 4424, 10556, 16832, 5364, 1324, 4504, 30990, 27290, 14412, 19356, 11134, 27132, 23222, 12468, 12060, 6782, 15840, 6550, 1638, 0, 13670, 36688, 27104, 35672, 14330, 1210, 21932, 25130, 31236, 25348, 26978, 18994, 20626, 33214, 30150, 32608, 30620, 32962, 29380, 36070, 14972, 1064, 25440, 19242, 14028, 16570, 15380, 18254, 14042, 26266, 20484, 16794, 25004, 26986, 18254, 0, 4378, 16470, 27348, 29530, 31084, 32226, 32922, 32780, 32932, 35080, 35988, 35336, 36650, 35578, 34732, 35856, 32240, 30664, 30942, 32174, 29846, 27656, 29000, 28570, 28532, 29022, 27886, 30362, 20990, 3422, 0, 3102, 11176, 20012, 28128, 30560, 32140, 31428, 30548, 27712, 23462, 23584, 25612, 28432, 20472, 0, 7542, 2528, 8478, 7576, 5322, 13204, 0, 17038, 14528, 23676, 25930, 7068, 14816, 11178, 7152, 1756, 11410, 19596, 20344, 19770, 19024, 19596, 18642, 20466, 17004, 23766, 5660, 9554, 9698, 3816, 10308, 0, 3108, 0, 8858, 5552, 2896, 2838, 5394, 11772, 26038, 24054, 5154, 2436, 4374, 7832, 0, 27282, 28170, 15036, 20182, 19182, 19128, 26316, 34390, 21052, 1764, 5362, 15344, 15972, 21012, 22140, 22612, 14182, 8138, 9858, 9088, 9308, 9584, 8692, 10896, 9934, 21500, 33024, 31142, 34276, 18272, 14580, 27348, 31578, 26524, 23150, 29348, 29666, 38480, 30454, 19246, 26308, 29414, 30212, 31422, 31330, 29846, 28022, 17468, 21244, 18660, 14164, 8526, 0, 13990, 10382, 0, 12638, 5562, 8268, 9222, 4054, 19430, 13820, 16118, 16038, 14008, 19006, 4866, 8020, 14436, 4168, 29042, 24490, 23294, 24074, 13946, 7436, 0, 6116, 12400, 13124, 5542, 0, 1724, 0, 7078, 6828, 0, 4440, 0, 12542, 13278, 0, 9904, 16016, 13968, 13206, 13684, 9314, 18298, 22138, 13840, 15382, 14040, 14900, 14242, 14378, 14584, 13994, 15160, 12808, 20512, 28398, 27854, 31462, 31226, 32104, 32348, 31452, 32416, 31840, 32640, 32856, 37340, 23174, 21484, 23186, 18612, 26322, 23594, 25194, 16572, 18822, 25530, 21068, 25582, 32210, 30928, 30160, 32634, 33972, 33862, 33072, 34714, 36792, 34318, 34000, 35226, 36266, 37218, 37014, 36928, 37320, 36450, 38396, 30462, 10820, 0, 4666, 6222, 50, 6058, 6022, 11150, 22242, 14822, 16522, 25106, 27338, 18248, 12382, 13352, 10406, 11776, 10044, 8438, 606, 5516, 26300, 29936, 34238, 16424, 0, 10398, 23578, 25002, 24484, 22926, 20378, 18046, 29990, 24374, 12214, 16136, 14016, 15364, 14298, 15484, 13496, 20690, 32012, 21476, 15390, 23800, 32562, 24984, 21772, 22654, 15530, 21180, 28606, 15700, 1546, 0, 9874, 24188, 25378, 26710, 27586, 28298, 29306, 30498, 33344, 33380, 32210, 33230, 34740, 33196, 33040, 34728, 26814, 26034, 25108, 33408, 37854, 26486, 17572, 12708, 14274, 13224, 14330, 12698, 15712, 6460, 0, 0, 6310, 22306, 24852, 20102, 17836, 21212, 25162, 24380, 26384, 21728, 23690, 15888, 3278, 2492, 1030, 4992, 0, 25174, 13412, 3678, 8336, 2182, 16092, 12580, 18420, 24094, 24970, 4134, 7274, 23884, 28460, 32672, 33690, 26418, 14460, 14210, 13644, 14310, 13200, 15298, 11288, 19352, 1914, 16738, 21098, 9548, 16140, 8994, 8554, 19178, 19540, 16088, 30250, 24894, 28024, 31954, 17734, 0, 6814, 19132, 33788, 22320, 23388, 25058, 15788, 21434, 19130, 22530, 34706, 18020, 0, 1788, 0, 2034, 2098, 0, 3108, 188, 14472, 28652, 24322, 26456, 25380, 25804, 25800, 25836, 29086, 23432, 12254, 27360, 33540, 31542, 34738, 34906, 29200, 27548, 30232, 31850, 23034, 10276, 16530, 20470, 23406, 26184, 22876, 19488, 18686, 20238, 11132, 27926, 19954, 23084, 12992, 7246, 8866, 8014, 10164, 6338, 15372, 0, 11180, 5428, 3846, 13816, 10316, 11768, 11740, 10354, 13818, 3694, 7112, 23892, 18038, 26150, 26694, 12104, 3110, 0, 3582, 6194, 18792, 9994, 9768, 24178, 3452, 1760, 0, 13284, 8290, 7774, 13186, 13186, 30, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 70, 0, 245, 0, 2120, 5548, 5564, 5968, 6223, 5396, 5518, 2346, 0, 288, 0, 81, 0, 16, 0, 0, 1, 0, 8, 0, 26, 0, 448, 681, 342, 470, 178, 22, 69, 0, 13, 0, 7, 0, 20, 0, 70, 0, 818, 3348, 5054, 6345, 7071, 7192, 7982, 4591, 343, 41, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 12, 0, 41, 0, 532, 2308, 2987, 3431, 3610, 3609, 4247, 5179, 5065, 5088, 5625, 5459, 5846, 6063, 6406, 6058, 5387, 3129, 387, 0, 0, 0, 0, 0, 0, 12, 0, 71, 0, 251, 0, 2074, 4942, 4334, 4197, 3911, 3929, 4237, 2923, 1092, 449, 0, 62, 0, 14, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 17, 0, 59, 0, 493, 1181, 1313, 2575, 3578, 3812, 4164, 4508, 4549, 4547, 4547, 4547, 4544, 4547, 4605, 5225, 6090, 7200, 6945, 6375, 7584, 8164, 8423, 8280, 8673, 9151, 10837, 7483, 4032, 4779, 4089, 3454, 2791, 2298, 1525, 1012, 649, 816, 602, 819, 795, 220, 0, 17, 0, 0, 11, 0, 52, 0, 459, 1216, 1162, 1228, 1167, 1244, 1121, 1353, 596, 0, 63, 0, 0, 150, 980, 3579, 5636, 6838, 8631, 9409, 9896, 10359, 10327, 10337, 10535, 8497, 7011, 5679, 4258, 5048, 7452, 8958, 8439, 7754, 7378, 8093, 9408, 10194, 10622, 11091, 10981, 11379, 11302, 11023, 11081, 10952, 10947, 10980, 10889, 11076, 10720, 11437, 9083, 6053, 3339, 108, 81, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 559, 4561, 7941, 9075, 9608, 9693, 10227, 10275, 10362, 10338, 10339, 10346, 10338, 10352, 10109, 8798, 8397, 3251, 0, 310, 0, 110, 0, 93, 0, 821, 3190, 4646, 5026, 4996, 6105, 6858, 6322, 6397, 4825, 3540, 3843, 4610, 4974, 4300, 1507, 0, 175, 0, 83, 0, 134, 0, 1059, 2880, 4069, 6912, 7859, 7659, 7743, 7726, 7668, 7823, 7623, 8417, 3263, 0, 381, 0, 109, 0, 18, 0, 662, 5528, 9093, 8996, 9584, 9774, 9746, 9998, 10846, 12186, 11312, 12328, 6179, 774, 2536, 1710, 2231, 2049, 2421, 2077, 2384, 1064, 0, 133, 0, 38, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 34, 0, 126, 0, 1078, 3212, 5506, 8197, 8217, 8045, 7861, 7140, 6443, 4688, 1304, 0, 699, 1279, 1845, 875, 0, 111, 0, 32, 0, 6, 0, 4, 0, 19, 0, 67, 0, 570, 1376, 1250, 2219, 3413, 4348, 5614, 6835, 6286, 5728, 5805, 5535, 5505, 5274, 5062, 5292, 5445, 5299, 5166, 4890, 5044, 4958, 4859, 4274, 2241, 399, 0, 24, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 62, 0, 216, 0, 2050, 6414, 7351, 8164, 8586, 9132, 9790, 9913, 10843, 11865, 12352, 13550, 13623, 14067, 15001, 14284, 13327, 12602, 12066, 12881, 13854, 13879, 13909, 13897, 13888, 13920, 13872, 13733, 11284, 8230, 7904, 7367, 7497, 7475, 8187, 10036, 10965, 11996, 13532, 15144, 15250, 15201, 15946, 16742, 16679, 17058, 17154, 14871, 13749, 8414, 1145, 0, 91, 0, 1070, 4941, 7726, 8703, 8779, 8468, 7898, 7502, 7377, 7558, 7318, 6946, 7053, 7021, 7001, 7086, 6880, 7629, 8570, 8450, 8163, 8190, 4017, 1539, 3410, 4349, 6583, 7523, 7985, 8349, 9023, 9491, 10094, 10821, 10678, 11163, 10789, 10485, 9607, 13033, 16702, 15620, 13239, 12130, 13149, 13382, 13666, 13933, 14476, 15067, 15679, 16080, 16124, 15929, 15339, 14850, 15161, 14697, 15504, 14047, 16934, 7490, 0, 930, 0, 266, 0, 53, 0, 0, 0, 0, 17, 0, 84, 0, 298, 0, 2567, 6833, 7309, 7847, 7705, 8830, 9178, 8811, 7418, 7918, 3198, 0, 382, 0, 109, 0, 22, 0, 0, 0, 0, 4, 0, 25, 0, 91, 0, 796, 2210, 3162, 5739, 7585, 7736, 7974, 8110, 8456, 9047, 8864, 7953, 7642, 8236, 8524, 8768, 8780, 8520, 8601, 8217, 6899, 2165, 0, 226, 0, 64, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 95, 0, 336, 0, 2866, 7516, 7903, 8555, 8099, 8209, 8305, 8476, 8059, 7137, 7098, 5271, 1062, 0, 17, 58, 0, 726, 2083, 5944, 8522, 7998, 5721, 2051, 1489, 1702, 1299, 2066, 518, 5701, 11593, 10111, 10327, 9634, 9714, 8993, 8049, 2700, 0, 293, 0, 31, 115, 0, 836, 0, 3010, 0, 20093, 22907, 580, 11180, 7393, 10561, 9724, 10523, 10198, 10110, 10139, 10145, 10047, 9715, 8895, 8228, 6663, 5954, 6424, 7564, 8527, 8265, 8339, 8402, 8161, 9100, 10167, 9795, 9607, 9954, 8928, 7450, 2583, 0, 290, 0, 82, 0, 16, 0, 2, 0, 9, 0, 30, 0, 573, 3044, 4322, 6062, 8327, 8829, 9419, 8248, 7710, 8622, 9618, 9370, 8777, 7923, 5765, 4667, 3942, 3756, 3732, 3793, 3663, 3914, 3415, 4986, 6235, 5889, 6739, 4995, 4551, 5146, 5616, 6741, 7385, 7891, 7777, 8214, 7883, 8109, 7815, 7682, 7565, 6922, 6361, 4719, 2982, 961, 120, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 13, 0, 42, 0, 407, 1159, 249, 2769, 6153, 8245, 4537, 0, 488, 0, 3088, 6218, 5806, 6843, 5978, 6178, 6277, 7035, 2889, 0, 351, 0, 115, 0, 84, 0, 707, 2857, 4575, 5885, 7556, 8253, 5950, 4872, 5264, 5054, 5240, 4999, 5389, 4636, 7034, 9409, 9159, 5746, 3093, 4476, 4520, 4384, 3283, 2999, 3203, 5046, 7141, 8568, 9555, 10365, 12314, 13814, 14214, 14253, 14117, 14121, 14218, 14056, 13913, 13694, 13181, 13274, 13292, 12386, 11917, 10593, 9878, 3553, 0, 402, 0, 115, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 33, 0, 126, 0, 1234, 2637, 3536, 4482, 4534, 4583, 3675, 3656, 3578, 3165, 3388, 3656, 4041, 4584, 4368, 4347, 4760, 4941, 4875, 4950, 4831, 5038, 4626, 6064, 8203, 8570, 9246, 9417, 9523, 10084, 9907, 9994, 9418, 9069, 5914, 1537, 1885, 3531, 4027, 5718, 6506, 6546, 5334, 4373, 2439, 0, 2051, 4187, 6946, 8438, 9719, 7963, 4491, 5395, 4167, 3004, 2969, 4053, 4051, 6212, 9831, 10284, 10333, 10214, 10421, 10048, 10792, 8329, 5830, 6781, 6367, 6512, 6382, 6399, 6309, 6394, 6459, 6840, 5334, 1812, 350, 2154, 4618, 5644, 6353, 6812, 7343, 7603, 7396, 7522, 7419, 7294, 7354, 7310, 5629, 1222, 0, 0, 3032, 7221, 8891, 9532, 9537, 3632, 0, 462, 0, 317, 0, 719, 0, 5751, 14132, 14210, 16577, 16679, 17509, 17467, 17343, 17319, 17038, 16262, 14129, 13197, 13549, 13776, 14025, 13614, 13617, 13840, 14035, 14142, 14623, 14962, 15486, 15897, 16012, 15764, 15787, 15255, 14713, 14153, 13997, 11946, 12476, 5233, 0, 638, 0, 206, 0, 148, 0, 372, 0, 3302, 8687, 6751, 10706, 13734, 11763, 10261, 10254, 9515, 10610, 4501, 0, 465, 0, 0, 1856, 8982, 13424, 15236, 15176, 15728, 11404, 7575, 8797, 8682, 9128, 8921, 9110, 8784, 8707, 8918, 8936, 9158, 9234, 9498, 9700, 9772, 9984, 10006, 10056, 9944, 10158, 9760, 10562, 7839, 4554, 5077, 4650, 4844, 4987, 5023, 6108, 7768, 9427, 8359, 8630, 3660, 0, 451, 0, 128, 0, 23, 0, 0, 0, 4, 0, 5, 199, 2138, 3401, 3692, 4174, 4271, 3944, 5173, 6903, 7122, 7757, 8055, 8221, 8258, 8220, 8293, 8157, 8405, 7912, 9507, 10997, 10509, 10838, 10857, 11071, 11334, 11370, 12428, 13855, 14536, 15083, 15547, 15147, 14750, 14853, 14663, 14374, 14134, 14020, 13462, 11140, 9758, 10378, 10313, 10461, 10699, 10564, 11223, 12512, 12851, 14781, 14142, 15963, 6728, 0, 822, 0, 256, 0, 152, 0, 369, 0, 2980, 6800, 6095, 6158, 5827, 4932, 4363, 1435, 99, 0, 4383, 10764, 9562, 10635, 9820, 9871, 10286, 10027, 10008, 10155, 10071, 10345, 10429, 10760, 10696, 11192, 11803, 11599, 11227, 10667, 10143, 9622, 8783, 8853, 8641, 11651, 8457, 4027, 5324, 4674, 4986, 4910, 4776, 5161, 4423, 8081, 11708, 11953, 8488, 5877, 6956, 6806, 6665, 6164, 5022, 3733, 4274, 4427, 5352, 5877, 6090, 5971, 5678, 4336, 1734, 514, 1144, 1466, 1359, 1251, 1151, 1115, 1042, 1088, 1084, 1125, 1078, 1215, 709, 150, 116, 0, 20, 0, 5, 0, 0, 0, 0, 42, 141, 891, 1280, 7663, 14407, 15096, 15939, 15641, 17057, 18091, 18104, 18424, 18624, 18346, 17122, 16307, 14651, 13179, 12382, 11190, 5110, 1816, 2467, 2344, 1136, 0, 145, 0, 31, 0, 0, 52, 0, 196, 0, 1576, 3588, 2942, 3319, 3027, 3337, 2845, 4551, 6625, 2122, 0, 210, 0, 65, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 68, 0, 250, 0, 2043, 5150, 7028, 8851, 8719, 7722, 6925, 3216, 0, 187, 0, 151, 2410, 4520, 4529, 4772, 4706, 4667, 4825, 4496, 5077, 2109, 0, 255, 0, 73, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 29, 0, 100, 0, 1021, 3434, 4164, 5607, 7255, 7802, 7826, 7994, 7900, 8072, 6121, 5212, 3651, 325, 25, 0, 9, 0, 0, 0, 0, 0, 29, 0, 68, 139, 3301, 5464, 5880, 7225, 7536, 7822, 7992, 8262, 8462, 8676, 8224, 8445, 6401, 5924, 2739, 0, 979, 1592, 1725, 1448, 1475, 1422, 1452, 1400, 1449, 1368, 1447, 597, 0, 72, 0, 20, 0, 4, 0, 0, 0, 2, 0, 7, 0, 23, 0, 801, 5144, 7633, 8249, 10144, 10335, 10798, 11285, 11540, 11723, 11965, 11967, 11657, 11788, 11584, 11532, 11223, 11026, 10937, 10801, 11008, 11262, 11412, 11456, 11571, 11623, 11639, 11580, 11551, 11806, 11617, 11430, 11590, 11657, 12002, 12315, 12324, 12333, 12331, 12324, 12344, 12270, 12082, 11617, 11109, 10782, 10675, 10640, 10798, 10809, 10502, 8674, 6422, 3919, 718, 0, 40, 0, 11, 0, 2, 0, 0, 0, 0, 0, 11, 0, 55, 0, 192, 0, 1974, 6915, 8560, 9349, 9684, 10013, 10205, 10077, 10146, 10082, 10167, 10021, 10303, 9480, 9017, 8184, 7174, 6397, 5590, 5335, 5081, 5856, 6495, 8518, 9692, 9832, 9927, 9717, 9810, 9884, 9995, 10131, 10017, 9819, 9593, 9819, 10027, 10345, 10242, 9725, 9988, 9828, 9371, 8603, 6464, 1725, 0, 160, 0, 45, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 74, 0, 260, 0, 2398, 7202, 8538, 10524, 11373, 11222, 11507, 11454, 11882, 12318, 11628, 12228, 11237, 15169, 18697, 18193, 18130, 18938, 15183, 11752, 12943, 12581, 12907, 12248, 12385, 11876, 11577, 11283, 11076, 11162, 11069, 11209, 10959, 11468, 9710, 6671, 4562, 8408, 14132, 14745, 16118, 15065, 16016, 6299, 0, 740, 0, 177, 0, 153, 2503, 4098, 5529, 7049, 6082, 2047, 0, 225, 0, 57, 0, 0, 47, 0, 200, 0, 1584, 3736, 4978, 7007, 7655, 8284, 8122, 8184, 8196, 8109, 8294, 7915, 9132, 10179, 9957, 10863, 10599, 10402, 10563, 10657, 10472, 10097, 9730, 9063, 8313, 8164, 7180, 5591, 1804, 0, 195, 0, 51, 0, 0, 16, 0, 79, 0, 835, 3257, 4251, 4838, 4326, 5260, 2366, 0, 291, 0, 203, 98, 150, 140, 118, 172, 66, 380, 609, 745, 944, 1413, 4134, 6470, 6239, 7238, 3280, 0, 2479, 6230, 2473, 0, 266, 0, 54, 65, 366, 415, 302, 304, 402, 0, 507, 0, 4003, 9607, 8661, 9676, 9150, 9184, 9536, 9740, 9608, 9804, 9845, 9649, 9826, 9536, 10054, 9112, 10983, 4858, 0, 603, 0, 168, 0, 19, 6, 0, 74, 0, 958, 4180, 5565, 6114, 7071, 7896, 8221, 8380, 8493, 8387, 8955, 9795, 10675, 11374, 11575, 12000, 12393, 11929, 10632, 9341, 9225, 9186, 9331, 10193, 11225, 11938, 12354, 12533, 12470, 12527, 12467, 12538, 12429, 12997, 14591, 12476, 13020, 5436, 0, 665, 0, 191, 0, 42, 0, 17, 0, 127, 255, 282, 355, 337, 500, 438, 472, 609, 349, 484, 267, 0, 36, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 58, 0, 212, 0, 1767, 4310, 4546, 4390, 4720, 2132, 0, 306, 0, 213, 0, 1489, 5285, 6419, 6758, 7509, 8625, 9732, 10049, 9963, 10030, 9956, 10052, 9859, 10930, 13546, 8117, 3724, 5103, 4406, 4579, 4417, 4060, 3319, 1262, 0, 317, 369, 1089, 2224, 2764, 2930, 2783, 2941, 2301, 1687, 1954, 1969, 1884, 1879, 1667, 1247, 1137, 1035, 1067, 641, 36, 9, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 46, 0, 155, 0, 1327, 3360, 3360, 0, 0, 19, 0, 93, 0, 320, 0, 3170, 10268, 12159, 11848, 10990, 7755, 13726, 17882, 16578, 15387, 12334, 13310, 12503, 11785, 6490, 6123, 3214, 0, 436, 0, 121, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 5, 0, 289, 2092, 3297, 2978, 2647, 2603, 1370, 1966, 2587, 10445, 17944, 18340, 20310, 20421, 22297, 25299, 26830, 28098, 29812, 30596, 30688, 31026, 30515, 29139, 23062, 19327, 20510, 19665, 20599, 19213, 21799, 13513, 5673, 8521, 9445, 6313, 9187, 5939, 0, 832, 0, 234, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 125, 0, 437, 0, 3453, 7530, 5383, 5530, 4461, 5393, 2520, 9067, 16453, 14444, 14973, 14677, 14681, 14980, 14278, 15755, 10804, 4887, 3793, 1840, 952, 0, 128, 0, 27, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 72, 0, 255, 0, 2034, 4549, 4053, 4458, 4077, 4198, 4223, 4050, 4419, 3650, 6383, 10522, 11119, 15111, 18711, 23096, 25340, 26759, 25375, 28798, 15529, 3235, 7961, 6870, 8658, 9643, 11377, 10304, 9870, 9308, 8535, 6960, 5280, 4421, 3823, 2956, 2479, 946, 0, 110, 0, 31, 0, 6, 0, 0, 0, 0, 5, 0, 25, 0, 86, 0, 719, 1718, 1370, 1724, 1905, 2260, 1902, 2459, 1153, 0, 0, 658, 2066, 3351, 5537, 5957, 7455, 6659, 6268, 7580, 8920, 6823, 5602, 7134, 7949, 8674, 7226, 7274, 7197, 7375, 7620, 7958, 8022, 6872, 4885, 2472, 450, 0, 28, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 318, 3528, 9925, 12338, 12240, 11741, 12699, 5254, 0, 1112, 1127, 3164, 1032, 0, 105, 0, 37, 0, 6, 0, 127, 1183, 2372, 3177, 3625, 4706, 6854, 7351, 6843, 6350, 6013, 6183, 5972, 6311, 5713, 6886, 3051, 0, 400, 0, 274, 442, 1651, 3121, 3641, 3477, 3034, 3636, 3015, 3793, 1917, 0, 252, 0, 71, 0, 14, 0, 3, 0, 10, 0, 72, 94, 0, 65, 0, 446, 1020, 1172, 1195, 2248, 2648, 2744, 3495, 3153, 3452, 3068, 3734, 1643, 0, 204, 0, 58, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 113, 0, 392, 0, 3230, 7718, 6612, 6830, 5300, 3309, 1327, 375, 85, 0, 5, 0, 0, 6, 0, 299, 1348, 1984, 1707, 1099, 261, 0, 23, 0, 6, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 22, 0, 84, 0, 549, 473, 0, 0, 809, 2581, 3561, 3786, 6053, 8688, 7122, 8499, 10132, 16384, 21708, 20806, 20152, 19253, 20218, 20295, 20328, 20143, 19895, 18969, 18193, 16194, 19809, 19644, 15283, 14694, 15307, 17496, 15206, 18451, 19790, 17064, 17602, 16862, 17910, 16173, 19523, 8633, 0, 1072, 0, 306, 0, 62, 0, 0, 0, 0, 0, 0, 16, 0, 118, 0, 450, 0, 4323, 9020, 16010, 25490, 26462, 28814, 29997, 29667, 28993, 28486, 28652, 28332, 28642, 28587, 27561, 27409, 26551, 26271, 25298, 24671, 24901, 24693, 24972, 24519, 25390, 22511, 19179, 19254, 18230, 18157, 18098, 17799, 17246, 18673, 14573, 15731, 4584, 5663, 19370, 5202, 0, 387, 0, 147, 0, 46, 0, 0, 0, 4, 0, 13, 0, 27, 0, 395, 1604, 136, 3956, 6914, 6798, 3120, 0, 404, 0, 110, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 40, 0, 181, 0, 920, 1198, 3719, 9337, 7498, 13143, 18143, 16040, 15771, 11090, 3997, 0, 121, 0, 32, 0, 3, 0, 0, 3, 0, 19, 0, 61, 0, 755, 2353, 2549, 3057, 1741, 600, 1146, 901, 1602, 4337, 5667, 5387, 5406, 5599, 5122, 6150, 2710, 0, 271, 0, 0, 626, 442, 829, 3267, 2580, 5204, 10160, 18554, 24991, 25200, 27095, 28159, 27824, 28274, 27442, 27503, 28356, 28660, 28613, 28188, 27603, 26587, 25021, 23365, 23610, 24294, 26123, 27164, 26481, 25840, 22704, 18828, 18731, 19262, 19150, 19129, 19287, 18922, 19727, 16905, 13080, 12213, 12059, 4508, 0, 514, 0, 144, 0, 30, 0, 0, 3, 0, 21, 0, 73, 0, 1133, 1068, 0, 176, 213, 49, 356, 1647, 2136, 2355, 2420, 2500, 1852, 766, 328, 314, 175, 0, 20, 0, 0, 32, 0, 130, 0, 839, 768, 0, 278, 0, 58, 0, 13, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 13, 0, 47, 0, 390, 925, 861, 1562, 2035, 2073, 2344, 2460, 2461, 2409, 2527, 2297, 2764, 1224, 0, 152, 0, 43, 0, 8, 0, 0, 0, 0, 0, 1, 0, 10, 0, 47, 0, 304, 483, 1651, 2689, 3033, 2927, 3410, 4063, 4312, 4406, 4366, 1794, 0, 217, 0, 60, 0, 12, 0, 0, 1, 0, 4, 0, 12, 0, 1105, 8580, 13942, 12044, 9260, 8175, 5187, 3436, 4118, 2827, 2288, 2297, 1839, 3427, 5450, 2714, 1278, 860, 22, 286, 0, 54, 0, 296, 297, 0, 45, 0, 12, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 42, 0, 207, 0, 729, 0, 6329, 16684, 16453, 14838, 13321, 17108, 19578, 21344, 22074, 22192, 22606, 22555, 22456, 22342, 24800, 26400, 24830, 26760, 22761, 19970, 23361, 24095, 24602, 24646, 24084, 23429, 21231, 19179, 18925, 16753, 15781, 15422, 15028, 15330, 14863, 15681, 14208, 17128, 7577, 0, 941, 0, 269, 0, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 51, 0, 206, 0, 1433, 2331, 3914, 5415, 7996, 14321, 18782, 21751, 22148, 22895, 24157, 24896, 25792, 26608, 26438, 26603, 26356, 26814, 25941, 27621, 23521, 25054, 14733, 3529, 8357, 6881, 7797, 7947, 9701, 8866, 7242, 6246, 7445, 3195, 0, 399, 0, 135, 129, 2061, 1378, 0, 138, 0, 48, 0, 62, 59, 0, 24, 0, 291, 546, 697, 905, 1187, 1072, 2944, 4537, 3870, 4561, 3542, 5272, 1895, 13100, 25722, 23179, 24832, 24809, 26151, 26816, 27111, 27530, 27741, 27482, 27728, 28102, 28442, 29684, 29906, 29546, 28800, 27295, 28966, 29265, 31969, 29402, 36824, 15521, 0, 0, 15081, 37254, 28609, 31490, 9701, 0, 560, 6670, 15875, 14918, 16015, 15611, 15891, 15662, 15945, 15502, 16440, 11913, 428, 8492, 19264, 18744, 19052, 16220, 15710, 10812, 2471, 2570, 3719, 13660, 24246, 25900, 26652, 29190, 18847, 9032, 11629, 10674, 11321, 10552, 8892, 7051, 7409, 3413, 0, 183, 0, 56, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 151, 0, 527, 0, 4227, 10309, 10672, 9147, 982, 5466, 11276, 15663, 20344, 22838, 26793, 27184, 27553, 26319, 25148, 22897, 19442, 16904, 11381, 7601, 7496, 6938, 7075, 7171, 6814, 7643, 4743, 1170, 1515, 1446, 688, 0, 84, 0, 20, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 85, 0, 305, 0, 4028, 7167, 7331, 9218, 8674, 6892, 1485, 7054, 12116, 10874, 11096, 11672, 9905, 16688, 24454, 15647, 10913, 7693, 5188, 3409, 185, 65, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 40, 0, 153, 0, 1305, 3901, 6334, 7382, 7524, 14090, 17279, 16612, 16702, 17053, 16010, 20007, 24772, 20083, 17557, 19209, 21857, 21968, 26521, 27663, 34157, 19228, 0, 19665, 30631, 13053, 11879, 10514, 10899, 8387, 6435, 6385, 4982, 3618, 2432, 822, 0, 89, 0, 24, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 89, 0, 281, 0, 8243, 16486, 16482, 18019, 18324, 19038, 18235, 16752, 16085, 14351, 11091, 8517, 9848, 9465, 4761, 3350, 4113, 3653, 3304, 3525, 3839, 3343, 3295, 3223, 3051, 3299, 2838, 1745, 764, 115, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 60, 0, 188, 0, 3041, 5843, 4313, 7999, 8412, 8229, 10136, 9944, 11267, 11579, 10237, 8724, 8140, 6394, 4622, 2130, 9031, 17527, 18761, 21798, 22602, 24669, 27661, 28497, 29053, 29404, 29521, 28896, 26191, 24660, 25258, 24625, 25576, 23948, 27136, 16494, 4182, 6356, 4001, 2389, 1084, 1389, 1353, 1260, 367, 0, 35, 0, 10, 0, 2, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 7, 238, 1882, 878, 4343, 8286, 7912, 8179, 9975, 11236, 15538, 19342, 18224, 18716, 18558, 18453, 18891, 17233, 15686, 16331, 11391, 8875, 10437, 9065, 9125, 8328, 7310, 6850, 6603, 6395, 5295, 4544, 3702, 3527, 3996, 1601, 0, 187, 0, 53, 0, 11, 0, 0, 0, 0, 0, 8, 0, 41, 0, 1040, 6993, 13538, 15439, 15441, 15358, 15611, 15091, 16074, 14091, 20722, 27654, 23722, 23221, 22350, 21842, 21622, 21065, 20996, 19696, 19125, 18636, 18723, 18172, 18263, 20870, 24471, 22398, 21606, 23023, 21325, 21361, 20965, 20290, 14463, 12221, 11490, 11928, 5007, 0, 610, 0, 170, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 16, 0, 176, 855, 3097, 5942, 7621, 3333, 0, 270, 0, 174, 0, 2684, 5860, 7127, 8358, 8454, 9016, 9643, 9685, 9107, 6766, 6358, 2614, 0, 318, 0, 90, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 75, 0, 266, 0, 2814, 10376, 14295, 16160, 17194, 14928, 12896, 11507, 13471, 9287, 10205, 19658, 20257, 24251, 23051, 24245, 9916, 0, 1547, 0, 637, 47, 316, 213, 229, 285, 163, 353, 0, 2212, 7917, 13262, 5656, 0, 678, 0, 197, 0, 42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 7, 0, 62, 177, 193, 244, 512, 2153, 2540, 5274, 6819, 9536, 12580, 11533, 12206, 11578, 12416, 10922, 15638, 20281, 17963, 11340, 6598, 6628, 2003, 14, 34, 0, 16, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 196, 0, 686, 0, 5540, 12442, 10462, 11225, 11224, 10464, 12438, 5548, 0, 714, 0, 431, 481, 557, 583, 452, 547, 398, 3019, 6156, 7823, 9587, 8110, 7587, 5714, 4066, 4968, 3062, 2681, 1903, 926, 552, 0, 83, 0, 20, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 20, 0, 97, 0, 396, 0, 1672, 2750, 496, 2093, 0, 4107, 13451, 15459, 20641, 24381, 25945, 27344, 26718, 27369, 26845, 25000, 24146, 20594, 17710, 7999, 0, 370, 0, 110, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 136, 0, 470, 0, 3898, 9390, 7981, 10053, 10638, 11553, 11093, 9258, 5571, 945, 22, 64, 547, 1037, 2353, 3288, 4376, 6067, 7922, 9283, 9966, 11092, 11262, 11352, 11126, 11559, 10757, 12377, 6697, 0, 1460, 785, 0, 91, 0, 33, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 107, 0, 365, 0, 3973, 14864, 17946, 17590, 18145, 18725, 18038, 2241, 7776, 19895, 16182, 17719, 17524, 16304, 21903, 27888, 25880, 25143, 21181, 16183, 8084, 3640, 1735, 221, 251, 0, 41, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 2, 0, 56, 0, 439, 602, 1984, 0, 8530, 20849, 23134, 26454, 25906, 26946, 27516, 24888, 22452, 22122, 20379, 15634, 4735, 0, 278, 0, 83, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 32, 0, 115, 0, 755, 772, 0, 156, 0, 354, 909, 750, 1002, 2037, 11200, 14652, 18444, 21177, 6008, 293, 1019, 2770, 7429, 9390, 8118, 6537, 7474, 6116, 5647, 4492, 1062, 0, 80, 0, 24, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 66, 0, 265, 0, 2150, 6258, 13096, 18068, 17068, 15655, 14230, 13212, 15039, 19554, 19652, 18144, 13470, 9351, 3598, 477, 1666, 1731, 2449, 3913, 6779, 7562, 7419, 7472, 7470, 7429, 7533, 7195, 7015, 7550, 7030, 7531, 2903, 0, 339, 0, 98, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10044, 11201, 8338, 18550, 30774, 29268, 30623, 30050, 30542, 30673, 31169, 31485, 31397, 31027, 30063, 28699, 29046, 30041, 29461, 27140, 23296, 17373, 14941, 10418, 5711, 3790, 8658, 14341, 16744, 19625, 19284, 19059, 20283, 24597, 26861, 27101, 27589, 28479, 28324, 28356, 28437, 28477, 28744, 28454, 28918, 28125, 29669, 24300, 17575, 20571, 12548, 7800, 8917, 6047, 9817, 15682, 18901, 19267, 20645, 19765, 22801, 26809, 26659, 27305, 27261, 28125, 28591, 28885, 29197, 29659, 29199, 28624, 29062, 26955, 22564, 20966, 16630, 13635, 14596, 9556, 5770, 6904, 4994, 11107, 18458, 18226, 18568, 18491, 18289, 18853, 17623, 21783, 26393, 25683, 26539, 27488, 28570, 28793, 26962, 26276, 25290, 22885, 23102, 18391, 14212, 14650, 9674, 5506, 5916, 4047, 7999, 15525, 16783, 17901, 18045, 18444, 20174, 23590, 26979, 27557, 28711, 28184, 29086, 29916, 29673, 30206, 30358, 29945, 29857, 29917, 30154, 29550, 30749, 28495, 33031, 18000, 2209, 7868, 11213, 16197, 16441, 18358, 18210, 18699, 21877, 22982, 22245, 23521, 23453, 24724, 25611, 24948, 25545, 26086, 26095, 25532, 23806, 22573, 22595, 17675, 14331, 15982, 10564, 5375, 6267, 4755, 7695, 12890, 13508, 15528, 15751, 16314, 19661, 20262, 20168, 20306, 20036, 20536, 19545, 22760, 25895, 25253, 25244, 24733, 22395, 20850, 19262, 16089, 14662, 14825, 8680, 4712, 6523, 4653, 10008, 14141, 14507, 16688, 16215, 18571, 20722, 22581, 23766, 22845, 25526, 26209, 25799, 26849, 25672, 25461, 25246, 22766, 19948, 19023, 17555, 16081, 15978, 15188, 15490, 15320, 15439, 15322, 15489, 15162, 15892, 16262, 15886, 18473, 21733, 23479, 23357, 23110, 23861, 24737, 24839, 25078, 26393, 24654, 22452, 19981, 18969, 18256, 17602, 16483, 15979, 9881, 6304, 9613, 9064, 7996, 11479, 15161, 15532, 16713, 15847, 15735, 17763, 20177, 20737, 21768, 22419, 22513, 22559, 22437, 22673, 22245, 23100, 20107, 16319, 17975, 14691, 9202, 6381, 5482, 5766, 6916, 6574, 8097, 12319, 14190, 15714, 15596, 14933, 14371, 15104, 16238, 15185, 17708, 20207, 22072, 20061, 16767, 17062, 16365, 17134, 16493, 17215, 15378, 11626, 7217, 4062, 4588, 3559, 6217, 6659, 5201, 5639, 5576, 5308, 6019, 4468, 9675, 15017, 13766, 14045, 14880, 15704, 15572, 16017, 15948, 16486, 16734, 16002, 16947, 13266, 9797, 7371, 3569, 4268, 3578, 3609, 3989, 6179, 6265, 9388, 10414, 12200, 13617, 10695, 12177, 12177, 12735, 13158, 14118, 15080, 15560, 15790, 15899, 16238, 16148, 16302, 16034, 16511, 15646, 17396, 11105, 1680, 3949, 5857, 5861, 5260, 6667, 9439, 12690, 12492, 10955, 11742, 11095, 12441, 13723, 13096, 14366, 15038, 15236, 16060, 15369, 16304, 13146, 9925, 10184, 7627, 5859, 5191, 5194, 3762, 3360, 2621, 4983, 3840, 3370, 6930, 9660, 11913, 10807, 11250, 11109, 11025, 11358, 10595, 13229, 16238, 15834, 15849, 15513, 12069, 8907, 7603, 6002, 5480, 4969, 4538, 4073, 3653, 3841, 5670, 5400, 6666, 8997, 10769, 11826, 11157, 11847, 13150, 13133, 15810, 15088, 13938, 15269, 15378, 15603, 16591, 12364, 8920, 8185, 5378, 5780, 4831, 4708, 4700, 4691, 4722, 4671, 4723, 5178, 9624, 12255, 12585, 15880, 17665, 17690, 18604, 17761, 17516, 15833, 15744, 16353, 15077, 17260, 16463, 13400, 7904, 5444, 6003, 5804, 5043, 5836, 7120, 6321, 7318, 10329, 11984, 12584, 12801, 15714, 19565, 18435, 17958, 18744, 18364, 18665, 17812, 16733, 17191, 16736, 17385, 16295, 18406, 11617, 5302, 7181, 6010, 5617, 6408, 8109, 5784, 10287, 13365, 13952, 14801, 16317, 19644, 19855, 19546, 19251, 19532, 19340, 18983, 18358, 17785, 18500, 19046, 19047, 19189, 17942, 18806, 13946, 7073, 6718, 6349, 7606, 9218, 6281, 10597, 15176, 14313, 15150, 14704, 15015, 14718, 15120, 14380, 16893, 20215, 19830, 19764, 19613, 19569, 20384, 20339, 20638, 18631, 18949, 11759, 4812, 6797, 6773, 9349, 7000, 8869, 14145, 15489, 15855, 16945, 17836, 18665, 19954, 20333, 20362, 20042, 20044, 20094, 20542, 20489, 21268, 20667, 21436, 21871, 19320, 18432, 18272, 18342, 18256, 18399, 18140, 18650, 16984, 15531, 16867, 16238, 16996, 17521, 18088, 20023, 20874, 21180, 20923, 19925, 20271, 20959, 20482, 21694, 21056, 20992, 22062, 19987, 17584, 18843, 10971, 4923, 6637, 7018, 9182, 7724, 12368, 16094, 15869, 17072, 17636, 18863, 19129, 20048, 21323, 21811, 21935, 21885, 21941, 21857, 22011, 21712, 22489, 21492, 18978, 18289, 17856, 10243, 5011, 7207, 8538, 8930, 9327, 14166, 16561, 16573, 17011, 18294, 18879, 19959, 21313, 21174, 22151, 21734, 21982, 21723, 21390, 20775, 21576, 22219, 21849, 21458, 19322, 17963, 18741, 11064, 4664, 7636, 8384, 9101, 8887, 9260, 8616, 9790, 7456, 14979, 21737, 19887, 22286, 21519, 22550, 22875, 22918, 21734, 21383, 22335, 22023, 22399, 21883, 19669, 17865, 19252, 11906, 5056, 7372, 9271, 8529, 11636, 16786, 16973, 17634, 17613, 18915, 20173, 20303, 20760, 22123, 23584, 22912, 22765, 23749, 23169, 22457, 22580, 22998, 22728, 23080, 22499, 23679, 18921, 8285, 7003, 9712, 9319, 10444, 15504, 17897, 17460, 17866, 18885, 19808, 20866, 21268, 21971, 22854, 22560, 22162, 22669, 22706, 22978, 22874, 22318, 22383, 22575, 21189, 19322, 18170, 19216, 10837, 5611, 9541, 8926, 9234, 14130, 18663, 17703, 18163, 18286, 18267, 18358, 18168, 18517, 17823, 20182, 23173, 22558, 23252, 23242, 23058, 22297, 22475, 22093, 20131, 18177, 19795, 11184, 5512, 9324, 9634, 7953, 12847, 19247, 17731, 18958, 18010, 18939, 19985, 20683, 21799, 23035, 23369, 22090, 22646, 22860, 22453, 23309, 24232, 24297, 23436, 23965, 21049, 18231, 18930, 18518, 18811, 18526, 18935, 17841, 17544, 18416, 18676, 18580, 19768, 21290, 21140, 22117, 22411, 23163, 22406, 22579, 23336, 24362, 24683, 23653, 23801, 23540, 23751, 22762, 19730, 19957, 15132, 8422, 9653, 9607, 10171, 15172, 18120, 18067, 18560, 18879, 20866, 21856, 22446, 23038, 23358, 23825, 23661, 23755, 23687, 23754, 23666, 23926, 24111, 23429, 23657, 21024, 19255, 17394, 10404, 8893, 10747, 9132, 14089, 19108, 17956, 19583, 19950, 20722, 21898, 22042, 23690, 24767, 24608, 24295, 24325, 24545, 24317, 23833, 24131, 23863, 23627, 23982, 23761, 23069, 22314, 21303, 15090, 10379, 10069, 9492, 9613, 9768, 9286, 10274, 8235, 15224, 23972, 23387, 24695, 24928, 24292, 24586, 24052, 23806, 24294, 23897, 24410, 24007, 24204, 24159, 21238, 19314, 18337, 9800, 7224, 10415, 9825, 12098, 16755, 19300, 19401, 19783, 20325, 20983, 23157, 23864, 23842, 24697, 24265, 23593, 23098, 22763, 23402, 24002, 23926, 23778, 24180, 23370, 25075, 18683, 7433, 7505, 9793, 10713, 11663, 16698, 19854, 19370, 19911, 19905, 20615, 22143, 23572, 23851, 24118, 23181, 22136, 21959, 21845, 22014, 22382, 23311, 23032, 22573, 20459, 18337, 19458, 14372, 8395, 8615, 9654, 9346, 14278, 19229, 18678, 18966, 19045, 19430, 19264, 19399, 19227, 19504, 18956, 20828, 23137, 22300, 21534, 21110, 21176, 22350, 23053, 21266, 21229, 20015, 20506, 13390, 8141, 8076, 10601, 17870, 17751, 20173, 22257, 22644, 20893, 20396, 21929, 22512, 23809, 24559, 24065, 24272, 25140, 23813, 22458, 21068, 19975, 21463, 21652, 20484, 20131, 19770, 19935, 19786, 19986, 19655, 20298, 18215, 16801, 19963, 22222, 20383, 20155, 22014, 23011, 24023, 22739, 23282, 24457, 24388, 22998, 22599, 21200, 20496, 23408, 22686, 21444, 20519, 19211, 15041, 9347, 7998, 8895, 7873, 12297, 17660, 16787, 18241, 20377, 19384, 18679, 20683, 21395, 22448, 22497, 21996, 22172, 22080, 22132, 22115, 22081, 22326, 22765, 21718, 17755, 18041, 12127, 7505, 9539, 8973, 7659, 12060, 17636, 16680, 17964, 19973, 19151, 19247, 21086, 22423, 22832, 23693, 25018, 24081, 24077, 22801, 21439, 22432, 23474, 24020, 22950, 21307, 18592, 17324, 10355, 5445, 7501, 6863, 6565, 5825, 5873, 6251, 5336, 7122, 3524, 15352, 27093, 23013, 25700, 24131, 23749, 23297, 21986, 21119, 21461, 22512, 22092, 22606, 19117, 18400, 9079, 1974, 5099, 5502, 3894, 7977, 15276, 15369, 18921, 20680, 20246, 22221, 23884, 24782, 24624, 24105, 24876, 25472, 25173, 24380, 23974, 23155, 23167, 22912, 23230, 22674, 23666, 21871, 25481, 12823, 0, 7737, 14631, 15728, 17200, 19851, 21061, 20887, 22681, 23157, 24146, 25025, 24382, 24806, 25930, 26536, 25916, 24920, 23840, 23390, 24307, 23839, 24139, 21776, 22317, 14021, 3523, 4303, 0, 7843, 16290, 15855, 19217, 21219, 21276, 22064, 23396, 22840, 23065, 22996, 22933, 23149, 22661, 24293, 25790, 24952, 24754, 25431, 25673, 25512, 23424, 22779, 12786, 4637, 3459, 9070, 17987, 19409, 21673, 21178, 23413, 23231, 22837, 23974, 24351, 25333, 27139, 26002, 25318, 26358, 25663, 25946, 25651, 23995, 24606, 26144, 25661, 26009, 22612, 21560, 14065, 7717, 9484, 8873, 8706, 9712, 7306, 15318, 22223, 20885, 24618, 23950, 25821, 27105, 26816, 26469, 27146, 27191, 26208, 26149, 25558, 25486, 26044, 25941, 25820, 23522, 20800, 15694, 8112, 13116, 18911, 18866, 21455, 21711, 22359, 22327, 21911, 23057, 23311, 23327, 25436, 26907, 26479, 26597, 26348, 25928, 26069, 25999, 26026, 26031, 26010, 25732, 23378, 22300, 19032, 12584, 15480, 20672, 21879, 23748, 24098, 23813, 22974, 22718, 24392, 24816, 24931, 25913, 26158, 27006, 27190, 26503, 27061, 27067, 27120, 27418, 26952, 27209, 26987, 26930, 25865, 23073, 22462, 17514, 15210, 20067, 22239, 22986, 23474, 23594, 23551, 23621, 23492, 23732, 23242, 25026, 27759, 26756, 26599, 27108, 26769, 26721, 27490, 27486, 28191, 28059, 27943, 25998, 22663, 23412, 18659, 13744, 17423, 20931, 21890, 22605, 22306, 22445, 21679, 20139, 20390, 21611, 22933, 23805, 23753, 24021, 24545, 24630, 24866, 25698, 25971, 26648, 27206, 26837, 27122, 26728, 27388, 26214, 28501, 21436, 17417, 22924, 21778, 22900, 22594, 21857, 21925, 22800, 23634, 24205, 25064, 25425, 25857, 25427, 25077, 25725, 26599, 27500, 27613, 27585, 27615, 25960, 25334, 23400, 21451, 17648, 11935, 13629, 16950, 19458, 22355, 22628, 23204, 23076, 21526, 22437, 23452, 23686, 23709, 23573, 23860, 23279, 25075, 26449, 27000, 27604, 26658, 26998, 26729, 25099, 24556, 20452, 17676, 13412, 6440, 12915, 18289, 18698, 20017, 19973, 20517, 20591, 20627, 21555, 22886, 23027, 22482, 23664, 24368, 24933, 26036, 25834, 26282, 25647, 25128, 24851, 24880, 22183, 20502, 19477, 17032, 17120, 17062, 16924, 17325, 16455, 19111, 20499, 20620, 21333, 21706, 23721, 24715, 24778, 24518, 26294, 26640, 26849, 26764, 27188, 25948, 25184, 25088, 25609, 22672, 20241, 19697, 17679, 15196, 8160, 6292, 8528, 14289, 18627, 19625, 20043, 19230, 20880, 22485, 24701, 26011, 26167, 26785, 27245, 27475, 27556, 27538, 27530, 27578, 27492, 27192, 22981, 20812, 19176, 17654, 12994, 7676, 7205, 10992, 16152, 18940, 21061, 20822, 20499, 21304, 22952, 23909, 24300, 24251, 25141, 25285, 25809, 26243, 26180, 26434, 24744, 23728, 23977, 23123, 19081, 17304, 17485, 17581, 10657, 5214, 8734, 8796, 14247, 18337, 17736, 18274, 17715, 18487, 17116, 21465, 25925, 25050, 25318, 25846, 26992, 26681, 26558, 25946, 25478, 25575, 25941, 23723, 18591, 17960, 15572, 8376, 6765, 8133, 9426, 13935, 18988, 20421, 20804, 19923, 21650, 23622, 23464, 24593, 25058, 25378, 26611, 26715, 26404, 26480, 26116, 26459, 26503, 26249, 26552, 25991, 27032, 25109, 28941, 16600, 5640, 10562, 13211, 18296, 19488, 20386, 19425, 21286, 22686, 23729, 24585, 25027, 25640, 25590, 26128, 27279, 26272, 25587, 25280, 25187, 25015, 24818, 20603, 16751, 19235, 15544, 10886, 9298, 8906, 9766, 13587, 19192, 20479, 20561, 20136, 21778, 23554, 23729, 23719, 23758, 23662, 23846, 23470, 24881, 27128, 25657, 25283, 25169, 23377, 19921, 17802, 19592, 15163, 7389, 7966, 10194, 10008, 14115, 18132, 18751, 18787, 19191, 21979, 23791, 24238, 25296, 26587, 27614, 27276, 27607, 28111, 27420, 26657, 26502, 26312, 26268, 24074, 20170, 17894, 19680, 14356, 9521, 10886, 10341, 10394, 10813, 9655, 13987, 20026, 20107, 22535, 24044, 25162, 25863, 25340, 25342, 25921, 26401, 26333, 25909, 26214, 25534, 25507, 23285, 19456, 17695, 19184, 12881, 7445, 9950, 10014, 10772, 14880, 18433, 17801, 18341, 18676, 22067, 24339, 25131, 26401, 26537, 26427, 25760, 26234, 26523, 26537, 26366, 26746, 26021, 27473, 22630, 17334, 17482, 9300, 7499, 10580, 10506, 10998, 15166, 18577, 18015, 18400, 18768, 21540, 23716, 24888, 26154, 26419, 26331, 26075, 26406, 26520, 26202, 26370, 26438, 25892, 24921, 20872, 17797, 18844, 15294, 7873, 8327, 11090, 10179, 12866, 17158, 18335, 18232, 18188, 18389, 17961, 18776, 17136, 22464, 27371, 25592, 27213, 26609, 26588, 26614, 25953, 25615, 23197, 20347, 17957, 18597, 14014, 6541, 8921, 10463, 10234, 14906, 18050, 17974, 18681, 17538, 19399, 23923, 25502, 26103, 26941, 26002, 25686, 26460, 26523, 26771, 26181, 26101, 24268, 22150, 20098, 18619, 19162, 18707, 19292, 18349, 20113, 14960, 13681, 18427, 17867, 18669, 18909, 20084, 23086, 26148, 26179, 26809, 26025, 25490, 26401, 26458, 26798, 26112, 25440, 23552, 22244, 20484, 18244, 16422, 9714, 6170, 8535, 9792, 9994, 11713, 16439, 18350, 18141, 17617, 18089, 21406, 24189, 26131, 26311, 26470, 26418, 26429, 26449, 26403, 26507, 26012, 24499, 23194, 20124, 18169, 16323, 9608, 6900, 8977, 9963, 10106, 14655, 18161, 17542, 17924, 19256, 20689, 23438, 24832, 25956, 27607, 27093, 27559, 27843, 27660, 28123, 27078, 25512, 26083, 24432, 22915, 19532, 17756, 14159, 7187, 8457, 10048, 9350, 9697, 9349, 9834, 9038, 10452, 7649, 16982, 27542, 26285, 27789, 27671, 28035, 27024, 28229, 28023, 26605, 26364, 26175, 25463, 23670, 19126, 19682, 12645, 6583, 10251, 9308, 9553, 15403, 18322, 19233, 21579, 21225, 23685, 24401, 25630, 27074, 27612, 27982, 27510, 27767, 28308, 28660, 26845, 25623, 25818, 25894, 25489, 26394, 24626, 28201, 16807, 7101, 9535, 12865, 18901, 19279, 22782, 21564, 22273, 23702, 24306, 25965, 27754, 28286, 28117, 28076, 27795, 27578, 28638, 28643, 26983, 26525, 26346, 25666, 23597, 19636, 20026, 12677, 7335, 10003, 9469, 14940, 20107, 21801, 21903, 21094, 22315, 23551, 23505, 23514, 23613, 23358, 23861, 22835, 26312, 30039, 27522, 26674, 26406, 26167, 24857, 22550, 18909, 18378, 12449, 8192, 10327, 9761, 15001, 20885, 22353, 23071, 23027, 23544, 23798, 25156, 26713, 27047, 27887, 27708, 27567, 27592, 28161, 28453, 27261, 26282, 26420, 25876, 24643, 19818, 18285, 16708, 14379, 15077, 14859, 14725, 15259, 14027, 18244, 22782, 22092, 24027, 24869, 26717, 27665, 28144, 27984, 27860, 28853, 28767, 28742, 27290, 26223, 26602, 26403, 25961, 20638, 18331, 16560, 8055, 7516, 7516, 0, 0, 0, 0, 0, 28, 0, 251, 0, 1023, 0, 5624, 205, 12761, 33638, 28498, 31018, 29931, 29874, 31077, 28338, 34033, 15180, 0, 2452, 280, 2084, 1856, 2636, 2880, 2433, 2725, 528, 2804, 0, 14675, 32593, 26191, 29318, 30405, 31484, 30409, 27158, 20727, 23207, 12986, 10729, 20753, 10700, 2657, 2374, 1137, 0, 122, 0, 36, 0, 8, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 81, 0, 603, 1029, 372, 176, 0, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 48, 0, 256, 0, 1163, 638, 14419, 28955, 29335, 26597, 22828, 24831, 24725, 27985, 24678, 33680, 17048, 0, 4932, 2608, 4618, 4216, 4813, 3936, 4493, 2419, 4614, 0, 14496, 31439, 24858, 27998, 27617, 28096, 27757, 28095, 27578, 28675, 23725, 9830, 3909, 3166, 2910, 1347, 0, 171, 0, 43, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 23, 0, 132, 199, 849, 1015, 73, 76, 0, 586, 1300, 1117, 602, 0, 33, 0, 9, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 250, 0, 906, 0, 4616, 971, 11169, 39477, 14501, 0, 1853, 0, 632, 0, 346, 0, 1394, 3556, 3485, 4161, 4451, 4861, 4583, 4125, 4015, 3730, 3691, 3657, 3823, 3425, 4065, 2364, 4256, 0, 12122, 25223, 18112, 20653, 16815, 14124, 5168, 176, 949, 0, 190, 0, 42, 0, 3, 0, 0, 0, 0, 0, 1, 0, 9, 0, 34, 0, 268, 695, 1248, 1514, 758, 162, 0, 20, 0, 62, 58, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 151, 0, 515, 0, 3807, 6714, 6090, 23740, 33116, 31460, 32802, 32229, 32511, 31856, 32215, 27008, 24360, 25132, 29266, 31108, 32659, 13082, 0, 3902, 2267, 4733, 3881, 4008, 3724, 3453, 2889, 3017, 2433, 3290, 1600, 4371, 0, 16676, 36846, 29972, 34568, 30041, 36676, 17143, 0, 4144, 248, 183, 0, 14, 0, 0, 16, 0, 43, 0, 162, 0, 965, 746, 1374, 4397, 3956, 5536, 7435, 9384, 12010, 9228, 5085, 3304, 783, 0, 153, 0, 20, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 30, 0, 257, 0, 1051, 0, 5366, 10, 13055, 34635, 29055, 34250, 29618, 36989, 16189, 0, 2490, 273, 3086, 2303, 2711, 2595, 2523, 2765, 2282, 3806, 4954, 4375, 4672, 4528, 3795, 4532, 2073, 4813, 0, 17156, 34098, 24906, 16928, 17146, 23628, 21930, 10195, 0, 1622, 0, 287, 0, 51, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 30, 2, 814, 1354, 1066, 1216, 469, 250, 246, 0, 40, 0, 10, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 137, 0, 455, 0, 9820, 25537, 28937, 32411, 29915, 36959, 16372, 0, 3579, 530, 2847, 1993, 2430, 2435, 2160, 2157, 2268, 1976, 3244, 4084, 4197, 4271, 3929, 4082, 3361, 4137, 2483, 4947, 0, 17025, 35560, 26199, 23906, 19276, 20354, 19080, 17315, 16087, 16516, 16125, 16669, 15767, 17506, 11946, 6965, 8972, 7867, 8551, 8740, 9317, 8391, 8733, 7142, 10816, 16800, 15750, 14159, 14943, 17481, 18465, 17093, 17024, 14717, 17922, 8479, 0, 1008, 0, 287, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 109, 0, 432, 0, 3211, 5007, 2079, 0, 9761, 27316, 29971, 31142, 32583, 28573, 35319, 16315, 0, 2863, 0, 1751, 1449, 2506, 3137, 3890, 4167, 4615, 4466, 4532, 4513, 4495, 4559, 4304, 4350, 3648, 3693, 1736, 4261, 0, 15088, 29980, 20074, 20393, 21497, 11241, 27, 3510, 1280, 1732, 978, 261, 0, 8, 0, 3, 0, 1, 0, 0, 26, 0, 140, 0, 500, 0, 3855, 8304, 8744, 10728, 8445, 8098, 8175, 7966, 8394, 7599, 9168, 4052, 0, 503, 0, 144, 0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 106, 0, 371, 0, 2956, 6853, 5383, 6643, 4998, 7654, 2632, 18003, 27778, 20486, 23470, 24809, 29904, 32840, 30603, 36352, 17347, 0, 4058, 1389, 2790, 2533, 1950, 3602, 0, 12009, 32248, 11815, 0, 4333, 0, 16634, 34783, 24872, 24131, 20892, 21471, 20762, 19914, 19238, 11860, 6402, 7042, 4948, 4391, 4153, 4275, 4139, 4362, 3960, 4771, 2110, 0, 261, 0, 73, 11, 485, 717, 877, 497, 1229, 822, 0, 110, 0, 9, 62, 85, 0, 12, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 213, 0, 904, 0, 4363, 0, 13920, 32463, 26282, 23651, 22661, 24192, 21413, 22134, 27065, 33155, 31582, 31040, 32191, 29692, 36892, 16110, 0, 0, 13110, 30753, 24526, 27215, 25838, 26371, 26468, 25772, 27357, 22974, 22043, 14068, 5528, 7346, 3511, 4662, 5058, 5083, 4751, 4229, 3974, 4023, 4452, 4476, 4254, 3812, 1254, 0, 134, 0, 38, 0, 54, 0, 234, 0, 837, 0, 6645, 14752, 12071, 4957, 0, 844, 57, 198, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 0, 401, 0, 1396, 0, 11908, 30593, 28634, 30116, 29256, 29729, 29457, 29719, 29248, 30723, 31686, 33025, 29566, 35811, 16793, 0, 4980, 3105, 4194, 3222, 3450, 3311, 2955, 3548, 1324, 4671, 0, 16359, 36161, 28151, 29381, 26823, 26145, 24577, 23664, 21285, 21360, 20497, 22396, 12310, 1139, 924, 0, 192, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 36, 0, 174, 0, 600, 0, 4388, 7048, 421, 229, 0, 315, 0, 3975, 19989, 27175, 25477, 25101, 25505, 9150, 0, 1026, 0, 291, 0, 51, 0, 0, 76, 0, 838, 1535, 2187, 2899, 2605, 2684, 2744, 2526, 3022, 1341, 0, 166, 0, 47, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 0, 438, 0, 1533, 0, 12658, 29992, 27823, 30688, 31827, 29301, 35764, 16387, 0, 3328, 88, 1898, 821, 1581, 748, 2961, 5083, 4268, 5134, 5043, 5036, 5103, 5240, 4600, 5216, 3460, 5350, 0, 16137, 37029, 28804, 30311, 28053, 27497, 23271, 21062, 17610, 11425, 9537, 4726, 121, 1534, 934, 0, 286, 0, 1218, 1108, 0, 36, 157, 0, 2021, 4636, 3824, 4255, 3968, 4223, 3909, 4339, 1756, 0, 209, 0, 60, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 60, 0, 286, 0, 937, 0, 8068, 21048, 13805, 8447, 0, 14042, 33140, 22956, 21360, 21207, 21363, 21325, 21519, 22306, 24403, 36884, 15697, 0, 3355, 0, 3545, 1716, 4910, 0, 15895, 28794, 31905, 17525, 0, 2612, 1997, 0, 16462, 35700, 26576, 22116, 16295, 17399, 16050, 16778, 16113, 17027, 15463, 18518, 8639, 0, 1721, 0, 427, 0, 81, 0, 2, 4, 0, 43, 0, 162, 0, 1247, 2902, 4138, 5134, 4095, 3228, 802, 0, 71, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 141, 0, 581, 0, 2893, 0, 8780, 26983, 28163, 28686, 29211, 26986, 33507, 14920, 0, 3887, 1025, 2555, 3088, 4901, 4469, 4714, 4624, 4654, 4671, 4552, 4887, 3856, 3776, 1733, 4967, 0, 16908, 32742, 19573, 22666, 20067, 22223, 13251, 5704, 7771, 2099, 0, 169, 0, 60, 0, 16, 0, 0, 0, 0, 0, 0, 0, 3, 0, 22, 0, 88, 0, 595, 1019, 2100, 3244, 2806, 3047, 2860, 3068, 2759, 3335, 1474, 0, 183, 0, 52, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 0, 556, 0, 1824, 0, 15188, 37527, 28709, 37492, 15229, 0, 4700, 1687, 4847, 4870, 5273, 5295, 5383, 5336, 5183, 5258, 4903, 4642, 4446, 3937, 4138, 3725, 4354, 2258, 4862, 0, 15925, 28794, 17363, 22648, 10973, 5347, 7079, 6718, 2615, 0, 306, 0, 78, 0, 16, 0, 0, 0, 0, 0, 0, 36, 0, 179, 0, 634, 0, 5045, 10856, 8491, 8158, 8301, 3551, 0, 286, 280, 931, 843, 601, 0, 82, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 140, 0, 516, 0, 11597, 14163, 4173, 0, 13671, 32881, 24280, 21964, 24640, 20652, 31629, 17094, 0, 4442, 1289, 2950, 3574, 4939, 4210, 4572, 4509, 4513, 4329, 4569, 4077, 5062, 3204, 6678, 0, 15859, 33294, 21394, 22314, 20446, 20110, 17728, 18986, 11844, 4110, 3634, 136, 110, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 189, 0, 808, 0, 3795, 0, 13429, 33698, 28921, 31642, 30045, 31128, 30109, 31656, 27051, 23967, 28014, 32148, 11994, 0, 3648, 1299, 2620, 2468, 2669, 1867, 1491, 243, 1701, 0, 2404, 0, 16114, 37242, 27677, 21766, 7297, 1756, 4182, 4929, 4975, 5026, 5373, 4795, 2886, 612, 0, 46, 0, 12, 0, 2, 0, 0, 0, 0, 1, 0, 2, 0, 126, 935, 1468, 1367, 468, 0, 52, 0, 14, 0, 1, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 38, 0, 123, 0, 1467, 4586, 932, 2618, 15219, 26592, 30022, 28842, 29989, 27778, 34374, 14432, 0, 5034, 1995, 3913, 3121, 3948, 3775, 3610, 2977, 2764, 2632, 2373, 2884, 3074, 2684, 1845, 2017, 1637, 1084, 1293, 1133, 1317, 1016, 1938, 2727, 1918, 1413, 1655, 747, 0, 92, 0, 25, 0, 5, 0, 0, 0, 0, 0, 26, 0, 137, 0, 475, 0, 3607, 7466, 6108, 8683, 4223, 2979, 2008, 0, 308, 0, 83, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 97, 0, 229, 0, 2251, 5150, 0, 14615, 26414, 18777, 22835, 20638, 22041, 21371, 21881, 21274, 22265, 20462, 24056, 12304, 764, 4747, 2371, 3596, 1125, 3533, 0, 17169, 35775, 24896, 33128, 12722, 1681, 0, 13908, 16561, 0, 5402, 2622, 6833, 7220, 7339, 7317, 7280, 7918, 6627, 5762, 2247, 0, 270, 0, 75, 0, 14, 0, 0, 0, 21, 0, 96, 0, 331, 0, 3019, 8357, 6831, 4245, 4145, 1847, 0, 228, 0, 64, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 152, 0, 592, 0, 3217, 3217, 30970, 28074, 33826, 14966, 0, 1870, 0, 588, 0, 312, 0, 1742, 4424, 4758, 4634, 5990, 7512, 7058, 7458, 7568, 7726, 7824, 7906, 7642, 7988, 7190, 8482, 3628, 0, 430, 0, 86, 0, 0, 746, 3190, 5410, 7282, 7454, 7034, 7546, 7790, 7770, 7710, 7868, 7546, 8182, 6384, 6618, 8670, 8042, 8628, 8744, 9184, 8880, 10412, 7806, 11474, 432, 12602, 28232, 23200, 29444, 27384, 30054, 30188, 30216, 30634, 30528, 30624, 29612, 29940, 30322, 26074, 27914, 31480, 30660, 31754, 32610, 32014, 31790, 31468, 31004, 31066, 31464, 31722, 31650, 31682, 31670, 31666, 31696, 31478, 30352, 28886, 28414, 29450, 31354, 31896, 31460, 32404, 31224, 30128, 27830, 28166, 26956, 24588, 25492, 26534, 28430, 28462, 28882, 29508, 26504, 31742, 12250, 0, 9070, 4930, 8598, 9248, 10070, 9480, 10576, 8114, 15694, 24762, 25074, 29510, 28420, 27404, 27658, 27548, 27564, 27654, 27380, 28406, 29822, 29666, 30864, 29814, 30218, 27130, 29066, 17596, 5046, 10112, 9618, 10906, 10168, 10620, 8960, 8910, 10902, 9828, 10586, 9488, 11382, 7516, 19320, 28680, 25150, 28386, 27530, 29738, 27966, 28984, 30470, 31210, 29990, 29074, 30280, 30024, 30612, 30562, 30602, 30600, 30570, 30632, 30516, 30882, 30808, 28980, 30080, 31440, 31532, 31456, 31952, 30454, 29192, 29484, 29152, 29822, 29312, 29672, 28672, 28336, 29726, 30710, 30224, 31666, 29034, 29846, 31572, 27086, 28682, 28430, 31402, 28676, 25356, 31254, 25642, 31966, 21882, 6552, 10544, 8670, 9654, 8864, 9182, 9082, 9062, 9176, 8940, 9722, 10422, 10076, 10268, 10074, 9714, 10408, 10224, 8584, 8666, 7534, 4852, 8120, 4056, 0, 682, 0, 732, 0, 4886, 12066, 11434, 12084, 9444, 10326, 11948, 11312, 11218, 10956, 10918, 10974, 10970, 10890, 11044, 10902, 10536, 10834, 10640, 10494, 10302, 10832, 9758, 11788, 7716, 20938, 33352, 29546, 31846, 30906, 31972, 32116, 31972, 31378, 28612, 27716, 19452, 3562, 0, 574, 0, 1386, 0, 11474, 29818, 24230, 26580, 15544, 6786, 10910, 8936, 12842, 9084, 18050, 14192, 20608, 32630, 25484, 29040, 28432, 30868, 33014, 33054, 31006, 31730, 31310, 31678, 31150, 32204, 29320, 29842, 26396, 35378, 9950, 10010, 11010, 4830, 10402, 0, 11484, 8536, 11394, 10906, 12332, 12084, 12196, 11774, 11332, 11422, 12264, 12266, 12150, 11012, 13438, 8472, 20830, 32674, 31126, 13092, 5074, 15178, 11466, 13360, 12544, 13314, 13474, 13780, 13514, 13634, 13536, 13650, 13478, 13808, 12542, 10324, 11698, 12894, 12812, 12810, 13270, 12672, 14398, 11862, 20644, 33142, 32322, 34106, 34142, 35500, 34426, 34458, 35232, 33962, 31034, 26978, 27996, 27338, 27042, 30744, 25802, 23626, 24656, 28606, 33382, 31954, 33866, 33376, 32542, 31744, 31814, 32278, 32090, 32236, 32070, 32312, 31900, 32976, 32248, 30118, 35140, 35126, 33760, 34942, 32996, 34492, 33378, 31840, 30080, 31114, 26926, 24352, 29050, 26262, 25366, 26008, 27334, 30034, 32940, 30312, 39880, 15760, 712, 14908, 10576, 14204, 13014, 15560, 11786, 23906, 37962, 35118, 34376, 33622, 33854, 34216, 35174, 35004, 34828, 35362, 34224, 37434, 36590, 32998, 37854, 34356, 35546, 34744, 38880, 26392, 12008, 17042, 14704, 16630, 16418, 17052, 16510, 15350, 16096, 17510, 15616, 17984, 12604, 26020, 39640, 34614, 36038, 34326, 34986, 35304, 34172, 27040, 32900, 30692, 30906, 37572, 33980, 33634, 27558, 28864, 31734, 30518, 31664, 30100, 32806, 25420, 25504, 32322, 33512, 33970, 34550, 38800, 37646, 39646, 40020, 40958, 38496, 37102, 37670, 36508, 35204, 37210, 28804, 30208, 28110, 20692, 26320, 26410, 27808, 31330, 33872, 30918, 29744, 23732, 22042, 27826, 32764, 29764, 35452, 13526, 1308, 14986, 13524, 17074, 15506, 16312, 15874, 16184, 15820, 16638, 15578, 13544, 14296, 13780, 14972, 16350, 15364, 16134, 12642, 11128, 11652, 15512, 7296, 0, 1182, 0, 1194, 0, 7842, 18946, 16386, 17756, 16452, 16706, 17458, 16330, 16070, 15968, 16104, 15574, 14768, 14854, 17622, 16246, 14906, 15168, 11020, 10274, 10004, 10734, 9296, 11994, 6568, 24504, 43020, 37580, 41100, 39756, 40408, 40582, 38702, 40136, 35254, 40594, 17988, 0, 2246, 0, 760, 0, 4146, 25254, 29376, 35124, 14578, 1738, 17404, 12964, 16512, 14238, 18284, 12872, 27024, 39622, 33206, 35862, 35944, 36906, 38898, 40428, 37526, 37102, 37144, 37032, 37282, 36810, 37798, 34564, 31888, 32344, 33838, 32176, 38368, 16166, 0, 1260, 2242, 12184, 13914, 15546, 15824, 16948, 17552, 17920, 17942, 17548, 19158, 19790, 20198, 19774, 16054, 16570, 13326, 27164, 41376, 37510, 38950, 32766, 40306, 16824, 0, 254, 6334, 19246, 15870, 16920, 16272, 16572, 16468, 16494, 16502, 16572, 17588, 18402, 18790, 18490, 19456, 18478, 19292, 20542, 22326, 17622, 30366, 44356, 39572, 40354, 38248, 39960, 38794, 38582, 38988, 38498, 28702, 25976, 28754, 26994, 34888, 25490, 22640, 24570, 26786, 33740, 32380, 38640, 39016, 35424, 36530, 35196, 37520, 40232, 39432, 39754, 39722, 39488, 40134, 37652, 34714, 38450, 36092, 36166, 37192, 29056, 28790, 27762, 25154, 22550, 20500, 23158, 21182, 16928, 16648, 21756, 21032, 25184, 25514, 26768, 36206, 30562, 39172, 14686, 3204, 20098, 15414, 19956, 18860, 20352, 18962, 21648, 17662, 33012, 44234, 37120, 40632, 39498, 40174, 39878, 39938, 40022, 39764, 40986, 43312, 38072, 35256, 38348, 39326, 42954, 39138, 43266, 27422, 13378, 20796, 18016, 20544, 21950, 21398, 20756, 21582, 22434, 19622, 24322, 39014, 45324, 42042, 41102, 39170, 37664, 35560, 35692, 38590, 37644, 37676, 35120, 36072, 37744, 33480, 25636, 29044, 33636, 32256, 32910, 32634, 32620, 32954, 31892, 31938, 30636, 34562, 39782, 36000, 39238, 42676, 42746, 42726, 41952, 40446, 40426, 40062, 38192, 35898, 33092, 33770, 34022, 33820, 30540, 31788, 38768, 31702, 34660, 37054, 32836, 33190, 22858, 25354, 25308, 29290, 34772, 42240, 18210, 0, 6298, 12776, 19326, 17204, 18110, 17888, 17568, 18542, 15822, 16994, 17436, 13630, 13904, 11078, 15628, 19534, 19962, 17518, 16390, 14800, 17318, 7262, 0, 0, 11534, 44698, 20306, 0, 10628, 20028, 18838, 18150, 16016, 16954, 18424, 16518, 16968, 16704, 16862, 15170, 12942, 17566, 19748, 16068, 14636, 13228, 12594, 12442, 13098, 11714, 14338, 9018, 27178, 47954, 37596, 39324, 43634, 41404, 40822, 40788, 41042, 42638, 40910, 39850, 39020, 36506, 35530, 31462, 30850, 29538, 28956, 37822, 33822, 42386, 16362, 2260, 18296, 16686, 16344, 26742, 41106, 38542, 40248, 40150, 40660, 40634, 42490, 41040, 42336, 41836, 40094, 40722, 40332, 40658, 40274, 40918, 38852, 36282, 36026, 37056, 37848, 40538, 38000, 42302, 18898, 0, 8846, 15638, 17472, 18142, 19284, 20494, 20782, 21476, 20466, 20398, 20780, 21060, 21846, 18964, 19884, 16274, 27626, 43868, 38762, 45324, 26596, 35306, 22096, 0, 1764, 4554, 20294, 19964, 20470, 20194, 20266, 20292, 20244, 20316, 20154, 20478, 21632, 22008, 21756, 22344, 21682, 21282, 22028, 25074, 19386, 33376, 45188, 40682, 42900, 42218, 45160, 42220, 42590, 39776, 38428, 29978, 30052, 27522, 27798, 29004, 17370, 20898, 21540, 25700, 32300, 34236, 38298, 40974, 39598, 40626, 38914, 40232, 42542, 41856, 42064, 42222, 41636, 42910, 39418, 40138, 40686, 34496, 41252, 38806, 38604, 32912, 26636, 28164, 25460, 35786, 23450, 17902, 17180, 15546, 23584, 21438, 26140, 23868, 34758, 37408, 43454, 18956, 0, 18280, 17054, 20882, 21504, 21536, 22388, 21730, 23050, 19420, 31392, 45576, 42092, 40124, 38232, 38792, 38686, 38448, 39076, 37748, 42026, 45180, 41232, 43558, 43134, 45102, 41654, 47334, 24820, 9676, 22432, 19072, 22170, 21246, 21524, 22440, 21604, 24510, 18086, 32490, 47092, 44526, 45054, 40708, 41062, 37138, 38214, 37772, 38652, 38684, 36442, 37348, 36810, 37244, 29778, 32572, 27712, 26250, 35172, 31936, 33582, 32698, 33218, 32832, 32494, 27524, 34662, 29022, 28108, 38138, 39064, 44034, 43058, 43556, 44026, 41426, 39262, 39894, 38444, 38522, 35022, 35992, 34262, 33628, 36650, 36494, 31070, 25928, 30212, 41838, 26394, 9980, 17702, 18368, 29674, 38540, 35862, 45510, 18638, 0, 1396, 5490, 14018, 11186, 12320, 12218, 11282, 15750, 22052, 17116, 13980, 13028, 14384, 18914, 19768, 17882, 16660, 11786, 18394, 6030, 16326, 58390, 12702, 18430, 47128, 44330, 19648, 2652, 25118, 18642, 17688, 13972, 16854, 16920, 17390, 16432, 15956, 15088, 13538, 14536, 20740, 17172, 11896, 12868, 12484, 15212, 15582, 16212, 14834, 17458, 12188, 29184, 43006, 33704, 41196, 44194, 42076, 39782, 40932, 41440, 43304, 38774, 44046, 19360, 0, 3970, 0, 14300, 32296, 34878, 36528, 43066, 20598, 0, 9626, 16370, 19430, 16848, 29284, 41504, 39388, 41842, 41710, 41660, 42322, 42450, 44790, 40432, 37908, 37554, 33920, 35284, 34518, 35042, 34524, 35822, 36880, 37456, 38718, 42496, 39144, 45844, 20336, 0, 6062, 12184, 18280, 17838, 19562, 20498, 21276, 21884, 21364, 21002, 21168, 22494, 21728, 19606, 20392, 15896, 27494, 41710, 41678, 41798, 38180, 40706, 36016, 18830, 0, 39508, 50968, 0, 2940, 0, 894, 184, 0, 1424, 0, 9870, 21582, 19166, 22214, 21256, 22076, 20444, 23212, 19310, 31448, 44364, 41922, 45402, 40652, 41010, 45780, 42372, 42556, 40242, 43982, 25876, 30570, 31344, 22344, 39708, 26602, 21312, 19850, 25872, 33732, 35316, 42158, 44682, 42810, 43592, 40786, 42458, 45684, 44200, 44956, 44426, 44946, 44218, 45542, 41602, 38434, 36228, 36598, 38122, 32566, 36744, 31474, 32012, 33044, 21932, 18034, 19686, 20914, 19072, 23078, 23232, 23640, 23728, 27552, 38624, 35508, 47540, 18978, 2172, 21764, 17564, 21636, 21186, 22310, 19776, 24562, 39296, 44422, 41742, 43884, 39732, 38830, 40972, 40128, 40680, 40188, 40764, 39832, 42674, 43746, 36898, 40048, 44878, 42842, 45310, 40276, 46064, 21450, 0, 13278, 22388, 21210, 21998, 21700, 22574, 20192, 26088, 41476, 44880, 45202, 42692, 41272, 40178, 37912, 39114, 39264, 38560, 36600, 36862, 36676, 37988, 39160, 32844, 34144, 35934, 30942, 30840, 30578, 30734, 30656, 30700, 30650, 30790, 31262, 34146, 38310, 40940, 41128, 42360, 42986, 42742, 44096, 41960, 38372, 37814, 39132, 36864, 34798, 35672, 35284, 35274, 35642, 30674, 27716, 35278, 37838, 35418, 37118, 18052, 12430, 18836, 23254, 32014, 31378, 31432, 41824, 17510, 0, 606, 8048, 19850, 15866, 17876, 16772, 17452, 16892, 17610, 14798, 12300, 13260, 12672, 17224, 19702, 18518, 15434, 14008, 8630, 0, 17526, 57116, 13270, 18654, 48404, 44558, 22944, 0, 3494, 11262, 22354, 18368, 20838, 20842, 17166, 13402, 15776, 14500, 13994, 13050, 16344, 16358, 12258, 13514, 13846, 16008, 16542, 16164, 16900, 15512, 18072, 12976, 29528, 45530, 41874, 44946, 44300, 42448, 39328, 41576, 43314, 40616, 37674, 36938, 36060, 35772, 33310, 31352, 25470, 28502, 35106, 36174, 35438, 33548, 8998, 4536, 18628, 14650, 18426, 31960, 39688, 38352, 40582, 39802, 40452, 41264, 43132, 41098, 38794, 36498, 34756, 35286, 35024, 35164, 35082, 35182, 35160, 36546, 35804, 39488, 38932, 41288, 26516, 1564, 878, 0, 7412, 16390, 15872, 16406, 18810, 19664, 19574, 17680, 15808, 19454, 17682, 18746, 15858, 21158, 2212, 18580, 48040, 40144, 42848, 39722, 37724, 42762, 17848, 0, 2142, 0, 614, 0, 184, 0, 284, 0, 994, 0, 8078, 18654, 16300, 18010, 17980, 17762, 21034, 16294, 29690, 42662, 37620, 41548, 40680, 41740, 43150, 40540, 38414, 36446, 35392, 37692, 32210, 31386, 24048, 24308, 39348, 27208, 15820, 23728, 27440, 35246, 26794, 32748, 42360, 35188, 37958, 36606, 39252, 41464, 42522, 42316, 42310, 42462, 42112, 42866, 40246, 37872, 41516, 39618, 30902, 32768, 38638, 36046, 24532, 18314, 30044, 35618, 34378, 24094, 21588, 29674, 23444, 28324, 30940, 36788, 38484, 43720, 19746, 0, 2142, 0, 0, 6454, 21338, 10718, 30694, 32378, 27098, 42824, 37152, 41398, 39446, 39750, 40726, 40396, 40502, 40602, 40242, 41062, 38306, 35834, 41072, 41538, 42516, 38506, 45264, 18858, 0, 294, 6922, 20584, 17612, 19392, 19082, 18422, 20114, 10828, 24736, 42476, 38792, 41878, 37496, 38162, 37186, 36862, 35036, 33972, 36210, 35674, 35606, 30314, 27974, 27364, 24594, 23674, 23896, 24724, 24790, 24758, 24858, 24642, 25064, 24220, 26746, 28394, 30556, 33834, 37394, 40456, 40548, 40862, 41858, 37806, 36196, 38734, 35146, 36354, 33000, 31818, 29210, 26308, 20360, 22484, 30142, 28192, 27412, 28582, 25712, 13770, 19386, 22266, 21416, 27090, 32748, 32158, 38112, 16860, 0, 2092, 0, 574, 0, 0, 242, 0, 1050, 0, 7884, 14754, 10982, 16534, 17412, 18406, 16240, 9278, 0, 21704, 47278, 41480, 44222, 40312, 42774, 37076, 45084, 18886, 0, 784, 5098, 17566, 16550, 17488, 17064, 14690, 12398, 12442, 12038, 11442, 13434, 13088, 11058, 10510, 11188, 15638, 14944, 12980, 12894, 12580, 13216, 12042, 14196, 9872, 24388, 41028, 37588, 36324, 34000, 33816, 38164, 38840, 33922, 34066, 33742, 33740, 31372, 29796, 27746, 27826, 30842, 36352, 32750, 36604, 14964, 0, 9944, 15204, 2094, 14098, 36368, 31950, 37782, 36094, 38366, 38208, 38056, 36490, 33282, 33774, 35548, 34558, 34370, 34372, 34354, 34414, 34346, 34392, 34494, 35716, 38854, 34408, 39154, 16276, 0, 1206, 2380, 11310, 11346, 12252, 12604, 12992, 14150, 11470, 8988, 12646, 14472, 13696, 14964, 8604, 0, 16262, 39764, 36320, 40742, 29460, 25770, 40286, 14934, 0, 1626, 0, 496, 0, 92, 0, 0, 242, 0, 840, 0, 6762, 15514, 12064, 14304, 12670, 15458, 10074, 23456, 37826, 33316, 36808, 36948, 37764, 39380, 36016, 33222, 33748, 32502, 33644, 23150, 19998, 17520, 26824, 27854, 17484, 20730, 20884, 22324, 27124, 31244, 31976, 35226, 33938, 35068, 33834, 37034, 39814, 39218, 39146, 37970, 38178, 38490, 37548, 39624, 33452, 32262, 34312, 34940, 30130, 28612, 27604, 18162, 27508, 29664, 27098, 27200, 27394, 26706, 23932, 21482, 25280, 29854, 31672, 35562, 34132, 43150, 17500, 0, 600, 1712, 0, 16702, 10368, 13026, 41746, 31644, 37836, 35074, 36674, 35636, 35020, 37330, 35708, 33320, 34164, 33572, 34188, 33250, 36138, 39134, 39248, 38312, 39492, 36086, 42060, 18582, 0, 3096, 0, 6470, 7704, 0, 938, 536, 22122, 37690, 34004, 35790, 35930, 37074, 35120, 32920, 30724, 32838, 27946, 29100, 33178, 32580, 28722, 28924, 29994, 24574, 26050, 21094, 21170, 21040, 18894, 19664, 19280, 19450, 19440, 19236, 20748, 28046, 36282, 38732, 38384, 39286, 39598, 38736, 37036, 36176, 36562, 33644, 33196, 29652, 24934, 26410, 22942, 18400, 18720, 28984, 28028, 20878, 21550, 29660, 29660, 21913, 21756, 23217, 23977, 25878, 27238, 28137, 29206, 29216, 29816, 29482, 28908, 28445, 28806, 28208, 29287, 27319, 31232, 18353, 4991, 8670, 6160, 8102, 7495, 6640, 5250, 4086, 4607, 3344, 824, 0, 68, 0, 18, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 26, 0, 94, 0, 625, 643, 0, 91, 0, 25, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 8, 0, 31, 0, 212, 169, 162, 353, 1010, 0, 2028, 1665, 8580, 14932, 10821, 14686, 20281, 35082, 16568, 0, 3157, 3223, 0, 14633, 32532, 26043, 29673, 27322, 28108, 26821, 26901, 27410, 27224, 27213, 27195, 27255, 26908, 26704, 26646, 26540, 26519, 26529, 26509, 26547, 26473, 26692, 26796, 26787, 26840, 26776, 27011, 27286, 27225, 27300, 27471, 27550, 27562, 27397, 27396, 27367, 27333, 26936, 26337, 25945, 25914, 26518, 26223, 26123, 26151, 25769, 26780, 24115, 20618, 18974, 17798, 13077, 2671, 0, 0, 2407, 6107, 4833, 5344, 4317, 3754, 3823, 3929, 3616, 4319, 1920, 0, 238, 0, 68, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 29, 0, 141, 0, 486, 0, 4285, 11577, 11336, 13205, 14002, 13736, 15244, 15838, 10930, 7835, 8199, 6499, 5787, 6341, 6181, 6189, 6178, 6723, 5854, 5581, 2292, 0, 240, 0, 0, 812, 0, 3160, 0, 23392, 15533, 10606, 38144, 22844, 20269, 15185, 6725, 0, 885, 0, 664, 0, 1628, 0, 12758, 28780, 23922, 25803, 23349, 23472, 23804, 22651, 21846, 21754, 24311, 26717, 29068, 34285, 30291, 36791, 15969, 0, 3173, 1239, 930, 2371, 0, 15002, 34394, 24039, 24156, 22996, 22489, 22514, 23147, 22305, 22719, 23589, 22902, 22525, 22460, 22743, 22636, 22738, 22587, 22853, 22369, 23327, 20534, 19920, 21352, 19957, 20356, 21990, 16408, 3201, 0, 196, 0, 60, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 0, 204, 0, 722, 0, 4795, 5140, 0, 663, 0, 219, 0, 203, 0, 613, 0, 5094, 14489, 19010, 27079, 25787, 33868, 15878, 0, 5185, 2452, 4233, 3419, 3401, 3075, 2544, 3177, 1644, 3632, 0, 14690, 31724, 26534, 29110, 27762, 28393, 28234, 27926, 28402, 28425, 26882, 27549, 28038, 28140, 28910, 29093, 29082, 29159, 29178, 29401, 29500, 29530, 29495, 29907, 29032, 30345, 27720, 35349, 18114, 0, 6776, 0, 16340, 35665, 26196, 27901, 21242, 17053, 17142, 16552, 16454, 15641, 14710, 15014, 14014, 12959, 13113, 13386, 12576, 14237, 10991, 19229, 10954, 0, 1485, 0, 422, 0, 83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 0, 94, 0, 309, 0, 6194, 19274, 23523, 29011, 28246, 34579, 16045, 0, 5589, 3148, 5176, 4366, 4811, 4761, 4898, 4877, 4833, 4585, 4592, 4615, 4496, 3485, 3185, 3128, 3709, 2443, 4871, 0, 16094, 32244, 27019, 29122, 27934, 28619, 28221, 28343, 28287, 27979, 27612, 27609, 27751, 27866, 27755, 27725, 27863, 28146, 28465, 28247, 28877, 28373, 27037, 27212, 27263, 27439, 27507, 27517, 27962, 27915, 28204, 26983, 25124, 24202, 23240, 21743, 17931, 16472, 16882, 16717, 16783, 16808, 16668, 17016, 15916, 14900, 13320, 13726, 9305, 4874, 8521, 6472, 4357, 5276, 5110, 5968, 2863, 0, 189, 0, 57, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 202, 0, 851, 0, 6346, 15681, 31054, 16848, 0, 4790, 1280, 3241, 2656, 3190, 3259, 3312, 3923, 3797, 4285, 2514, 5082, 0, 16395, 34540, 29026, 31709, 30404, 30825, 31181, 28889, 26173, 27096, 26818, 26477, 26693, 26813, 26977, 27524, 27287, 27442, 27728, 27675, 27778, 27677, 27785, 27831, 27961, 28330, 28485, 28868, 29027, 29366, 29168, 29064, 29060, 28989, 28698, 28754, 28846, 29035, 29300, 29370, 29493, 27102, 24150, 21229, 16069, 13785, 14514, 13879, 14728, 13350, 15992, 7261, 0, 2106, 2025, 2296, 2500, 2703, 3008, 2312, 771, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 73, 0, 263, 0, 2494, 7283, 7693, 8979, 15809, 21866, 24589, 26884, 26879, 27338, 28403, 27902, 30562, 27850, 34941, 15965, 0, 1234, 1290, 0, 14243, 33190, 27450, 29523, 27876, 29018, 28558, 28816, 28723, 28744, 28739, 28730, 28757, 28671, 28599, 28584, 28569, 28687, 28731, 28847, 28863, 28983, 28995, 29074, 29119, 28647, 28262, 28218, 28327, 28273, 28153, 27767, 27490, 27346, 27003, 26790, 26469, 27371, 25497, 26672, 10344, 0, 1212, 0, 348, 0, 71, 0, 0, 0, 0, 33, 0, 167, 0, 579, 0, 4655, 10676, 9117, 11354, 9142, 8716, 7810, 6966, 3010, 0, 378, 0, 103, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 0, 278, 0, 1043, 0, 8424, 19329, 23443, 27047, 34777, 16117, 0, 4373, 1673, 3727, 2847, 3045, 2800, 2593, 3239, 1958, 4355, 0, 15352, 31417, 26870, 29305, 28031, 28620, 28280, 28367, 28215, 28072, 28103, 27980, 27831, 27851, 27845, 28024, 28140, 28123, 28150, 28542, 28625, 28526, 29075, 28420, 29742, 27821, 31196, 17464, 2305, 2475, 0, 466, 0, 102, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 170, 0, 888, 0, 3158, 0, 20665, 20565, 0, 3705, 0, 1379, 0, 765, 291, 85, 0, 0, 62, 0, 320, 0, 1116, 0, 9232, 22126, 19426, 23099, 24259, 25197, 25868, 25776, 26599, 26359, 25404, 25555, 25491, 25456, 25605, 25259, 26414, 27483, 27321, 27936, 27930, 27802, 27549, 27384, 27159, 26872, 26505, 25867, 25726, 25816, 25922, 26028, 26151, 25766, 25718, 26762, 27322, 28014, 28128, 28159, 28366, 28618, 28640, 28390, 28236, 28541, 28842, 28929, 28656, 28809, 27242, 24165, 23109, 22605, 22507, 22611, 22399, 22801, 22078, 23508, 18648, 12612, 14112, 10786, 9799, 3930, 0, 481, 0, 137, 0, 26, 0, 0, 0, 2, 0, 10, 0, 83, 164, 261, 143, 0, 19, 0, 5, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 141, 0, 371, 0, 6596, 20956, 21911, 31462, 14769, 0, 3856, 2551, 4719, 4138, 4175, 4825, 3393, 5762, 0, 16017, 31871, 26121, 28809, 27401, 28168, 27758, 28007, 27770, 28153, 26875, 25402, 25578, 24934, 25584, 26215, 26341, 26568, 26529, 26686, 26952, 27066, 27132, 27330, 27534, 27715, 27705, 27746, 27416, 27503, 27853, 27950, 27970, 27868, 27729, 27947, 27853, 27822, 27490, 28151, 27702, 28449, 25963, 30381, 13205, 0, 1628, 0, 471, 0, 124, 0, 105, 0, 1223, 4813, 6319, 6714, 7219, 4382, 2628, 3531, 3468, 3006, 4277, 2068, 0, 262, 0, 75, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16301, 14527, 14747, 14797, 14545, 13598, 14032, 14253, 14785, 14696, 15824, 10951, 5370, 4394, 8363, 12174, 11031, 11547, 11356, 11309, 11623, 10649, 11359, 12046, 9587, 13806, 21165, 14314, 7695, 9209, 7708, 7468, 7284, 7603, 6980, 10861, 12650, 13865, 12960, 8654, 8329, 4758, 3383, 1364, 0, 195, 0, 146, 0, 350, 0, 3166, 9037, 9339, 13169, 18147, 10206, 3015, 5810, 6163, 6406, 6009, 6668, 5397, 9383, 12460, 11621, 13979, 13644, 14702, 14358, 14037, 13944, 15517, 16098, 15930, 16433, 15154, 13849, 11852, 8102, 5177, 5310, 5532, 6881, 7533, 7564, 7646, 7201, 6832, 7438, 7579, 5465, 6216, 2786, 0, 300, 0, 0, 267, 0, 2829, 8020, 7911, 8392, 7784, 8718, 6919, 13415, 24488, 26414, 27247, 27682, 26946, 28050, 26009, 22133, 21232, 20920, 16680, 14175, 14567, 14371, 14877, 14572, 15504, 15249, 14270, 12584, 12107, 10348, 8552, 6682, 5199, 4762, 4002, 3109, 2509, 2891, 2744, 3690, 4857, 4033, 5066, 9267, 1532, 6690, 16005, 12860, 14708, 13258, 14924, 11010, 9503, 9635, 6451, 6675, 8738, 6206, 15553, 25878, 25458, 26442, 24532, 24387, 23918, 22516, 21758, 20383, 23025, 17067, 11627, 15652, 15030, 15197, 14470, 14310, 12225, 9955, 7522, 6510, 5947, 5334, 4663, 4324, 3717, 3001, 2865, 2492, 2555, 2419, 2391, 2529, 2228, 2806, 1644, 5473, 9333, 7988, 8812, 9092, 8938, 7562, 5662, 7490, 8452, 8636, 7618, 13631, 19838, 18966, 19133, 17788, 18214, 18597, 18466, 18236, 18453, 19809, 17589, 13795, 13472, 14447, 16003, 15624, 13009, 10166, 6509, 3718, 4337, 4206, 4163, 4173, 3719, 3816, 3759, 3783, 3785, 3762, 3816, 3570, 2888, 2610, 2359, 3871, 5452, 4926, 6432, 8062, 7449, 8457, 8306, 7560, 7814, 7883, 7992, 7959, 6871, 9607, 14480, 17353, 18007, 16790, 17413, 12274, 9231, 10047, 11257, 12676, 12311, 11662, 9082, 6810, 6900, 8963, 9194, 6572, 4815, 4920, 4837, 4852, 4911, 4753, 5079, 4234, 4748, 4948, 3859, 4331, 3841, 4312, 5126, 4212, 3655, 4446, 4056, 3590, 3961, 2729, 4130, 6242, 5806, 7507, 9045, 8555, 8553, 6736, 11181, 17648, 13279, 8645, 12637, 10842, 10926, 12019, 8464, 6622, 1970, 784, 1364, 0, 1840, 4378, 3512, 4087, 3524, 4291, 2951, 6848, 8491, 5994, 6799, 5720, 6230, 6840, 6731, 6869, 6934, 6545, 5511, 4850, 6004, 5435, 4886, 5580, 5682, 6416, 4965, 6675, 6974, 3755, 6305, 7360, 7130, 6354, 6675, 3287, 452, 398, 215, 0, 3773, 8860, 5819, 13685, 12295, 6689, 8588, 7554, 8205, 7709, 8270, 6660, 3976, 3161, 2302, 6610, 9627, 6807, 6294, 7482, 7361, 9812, 11098, 11003, 10544, 8780, 8026, 6134, 6371, 6181, 5211, 5956, 3851, 2674, 2468, 3011, 4283, 4307, 4108, 4625, 3329, 7081, 6249, 186, 435, 0, 105, 0, 0, 67, 0, 377, 0, 1329, 0, 9362, 13825, 4947, 8209, 4539, 3995, 4417, 8338, 7345, 10037, 6949, 4936, 10296, 10337, 13188, 11682, 9633, 8984, 10492, 11802, 14099, 15110, 13036, 12957, 12718, 10600, 8294, 6534, 5536, 5361, 6335, 6014, 5357, 5422, 4182, 2479, 1058, 2484, 3335, 3147, 3168, 3291, 2962, 3690, 1423, 0, 0, 5050, 9451, 8924, 8315, 5225, 8201, 6558, 11167, 21536, 24343, 25004, 25450, 25388, 24743, 21153, 17257, 15597, 11913, 11473, 13074, 14143, 15246, 14819, 15019, 16217, 15786, 15833, 14310, 13349, 12323, 7925, 5949, 5310, 4653, 4800, 4689, 4731, 4733, 4703, 4761, 4627, 5481, 7896, 2979, 0, 88, 275, 0, 3954, 10256, 8621, 11095, 10710, 8482, 7880, 9182, 9553, 13655, 18866, 20111, 22388, 20430, 18818, 18943, 17758, 16866, 14352, 15630, 14183, 11251, 14256, 16940, 16842, 15805, 15833, 12634, 11314, 10238, 8467, 8467, 8410, 8384, 8517, 8236, 8809, 6911, 4978, 6057, 5251, 4709, 2421, 2391, 5361, 6619, 8002, 8295, 8739, 9392, 9469, 8541, 7860, 7099, 8531, 8626, 9350, 9447, 14013, 20461, 18905, 21343, 15874, 15823, 18232, 14111, 14718, 13680, 14556, 15014, 14986, 15099, 13891, 14632, 14482, 13391, 13860, 13450, 13975, 13138, 14731, 9563, 4357, 6167, 5451, 6354, 6792, 7245, 6249, 5415, 5162, 4731, 4021, 4785, 6108, 6125, 6182, 6361, 7674, 8192, 8260, 8326, 8677, 9102, 9080, 8667, 7907, 8695, 9414, 12648, 18130, 14249, 9659, 12738, 18242, 13642, 8759, 9693, 9423, 10646, 10200, 10368, 10387, 10186, 10673, 8941, 6451, 5771, 4309, 4830, 4768, 4413, 4969, 5069, 5631, 5873, 6317, 5827, 5747, 5201, 5564, 6106, 4927, 5067, 5679, 5290, 6181, 5723, 5055, 6520, 6744, 7161, 7160, 8116, 10354, 8147, 8369, 6929, 13288, 13289, 6305, 8383, 7235, 7893, 7640, 7616, 7901, 7270, 8556, 4530, 1783, 3917, 4889, 5468, 4220, 4770, 5887, 6946, 6932, 7605, 6880, 5607, 5660, 5645, 5546, 6495, 6801, 6850, 7101, 7278, 6503, 6956, 8126, 6748, 6342, 6753, 6870, 6706, 7340, 7797, 7755, 8197, 8326, 8372, 7678, 7249, 6416, 5853, 5946, 6040, 5731, 6373, 5086, 8809, 8853, 4518, 5442, 4605, 4335, 3526, 5492, 5129, 8333, 8543, 4470, 5335, 4641, 5258, 5452, 6219, 6758, 8438, 10047, 9814, 10128, 8983, 8072, 8312, 7808, 6783, 7103, 7036, 6343, 5848, 5514, 4801, 6069, 7756, 7575, 7852, 7927, 7958, 8037, 7830, 8241, 7474, 9001, 3988, 0, 503, 0, 163, 0, 933, 5942, 8029, 6999, 7471, 6244, 5527, 4508, 4511, 5488, 6146, 6553, 7768, 6077, 3090, 7276, 10116, 10657, 11980, 10476, 8845, 9362, 9663, 9824, 10240, 11378, 11548, 10285, 9348, 7955, 7170, 6416, 6100, 6163, 6163, 6109, 6283, 5270, 1876, 2220, 5291, 3907, 696, 0, 0, 118, 0, 467, 0, 3972, 9837, 8276, 9575, 8127, 7998, 9878, 7222, 9609, 10989, 18824, 28456, 28730, 28320, 26191, 24602, 24379, 18740, 16691, 13917, 10185, 12723, 12746, 13805, 13037, 13868, 14708, 14847, 14644, 15079, 14235, 15948, 10294, 4365, 5302, 4707, 5024, 4860, 5654, 6068, 5457, 5067, 5761, 5975, 7867, 4639, 0, 364, 0, 2372, 7039, 8094, 8721, 8925, 9399, 8675, 9115, 8932, 10063, 12113, 14422, 21134, 23887, 23413, 23050, 22309, 17488, 15503, 14049, 10259, 11297, 11554, 11539, 11584, 11484, 11689, 11011, 9717, 8159, 8265, 8072, 6766, 6470, 5861, 6185, 5808, 5412, 5234, 5219, 5051, 5413, 3058, 1376, 3787, 6162, 7720, 8030, 8532, 8140, 8911, 8786, 8052, 8494, 8171, 9518, 10287, 10677, 10284, 13039, 17648, 20040, 16703, 13727, 15127, 15341, 16100, 15759, 16028, 15705, 16256, 14508, 12521, 12215, 11058, 9795, 8313, 7263, 6982, 6890, 6924, 7200, 7032, 7088, 6386, 7084, 7561, 7123, 6587, 6048, 6231, 5865, 5421, 5708, 5487, 4617, 6005, 6244, 6803, 8363, 8358, 9594, 9767, 10028, 10619, 10141, 9143, 9610, 10890, 10834, 10936, 10835, 10977, 10734, 11195, 9995, 10780, 12605, 13427, 11518, 7270, 8448, 8593, 8352, 9053, 9204, 8029, 6603, 6491, 6326, 6560, 6702, 6601, 6524, 6647, 6615, 6490, 6467, 6667, 6624, 6718, 6248, 6149, 6721, 6559, 6775, 5907, 4781, 5060, 4883, 5606, 6370, 6608, 6859, 6750, 6848, 6719, 6932, 6517, 7834, 8880, 8313, 7028, 6855, 7013, 8623, 8398, 6635, 6033, 4386, 4472, 4380, 4994, 5538, 4728, 5208, 6374, 7446, 7851, 6912, 6574, 6168, 6202, 6172, 6279, 6539, 6540, 6823, 7499, 7356, 7490, 7438, 7096, 7457, 7541, 7491, 7495, 7507, 7534, 7459, 7620, 7300, 7930, 6259, 6195, 3133, 0, 163, 661, 3521, 4872, 8948, 8367, 5119, 5029, 4248, 4550, 4721, 5705, 6017, 6394, 7081, 7061, 6188, 5274, 5914, 6069, 6069, 7077, 7666, 7787, 8759, 9611, 9526, 9402, 9103, 7882, 6979, 7299, 7157, 7135, 7456, 7338, 7404, 7361, 7400, 7351, 7519, 7900, 7885, 7812, 7810, 7835, 4577, 551, 0, 0, 43, 0, 168, 0, 1749, 6161, 8570, 7290, 6906, 6376, 4894, 4965, 4404, 5192, 5707, 6910, 5821, 8506, 7022, 3855, 6198, 7539, 9791, 8234, 7598, 8606, 8500, 8263, 8055, 8156, 8040, 8220, 7909, 8520, 6459, 4158, 5769, 6033, 6607, 5272, 4823, 5581, 4279, 4064, 4142, 3823, 1187, 0, 87, 0, 0, 198, 0, 2116, 6889, 7778, 8767, 8538, 9466, 9208, 7542, 6154, 7480, 12211, 19581, 24483, 23740, 22674, 21637, 21087, 16920, 13276, 12854, 12882, 12824, 12967, 12676, 13270, 11464, 10017, 8077, 6426, 5917, 5553, 5939, 5460, 5730, 5002, 4285, 4348, 5047, 5826, 5596, 5782, 5561, 4109, 2698, 3984, 6762, 1660, 1431, 6575, 7635, 7824, 8806, 9374, 10281, 10174, 8309, 9568, 8763, 9874, 8425, 16043, 24278, 22054, 22760, 22424, 22364, 22850, 21775, 23989, 16827, 10259, 12181, 10707, 12266, 10241, 9660, 7711, 4993, 5382, 5097, 5687, 5705, 4446, 5354, 5841, 5528, 5433, 5264, 4628, 3889, 4608, 2691, 2207, 1587, 3694, 6934, 7919, 8390, 7637, 8099, 7944, 8406, 8316, 8700, 9530, 9948, 10193, 10232, 10175, 10301, 10058, 10507, 9613, 12560, 15467, 13834, 14166, 13716, 13365, 12415, 11743, 10339, 9185, 8986, 7512, 6847, 6901, 6498, 6066, 6185, 6467, 5498, 4489, 5557, 6168, 5138, 4544, 4947, 4915, 4201, 4186, 4436, 3829, 4636, 4611, 4719, 3868, 4707, 7905, 8189, 8222, 8220, 8191, 8267, 8120, 8389, 7863, 9542, 11086, 10637, 11069, 11060, 11802, 9875, 7243, 9000, 10080, 9311, 8524, 7815, 6728, 6655, 7954, 7746, 7146, 6734, 6274, 5301, 4957, 5148, 5173, 4907, 4696, 4640, 4703, 4536, 4540, 4961, 5065, 4972, 4021, 5142, 5669, 5077, 5150, 4757, 4908, 4838, 4861, 4872, 4823, 5009, 5237, 5257, 5952, 6477, 6345, 5632, 5251, 5018, 4418, 5063, 5692, 6203, 5245, 4983, 5193, 4850, 4511, 4122, 4228, 4711, 4474, 4565, 6078, 5606, 5608, 5748, 5238, 5164, 4924, 5021, 4833, 4896, 5041, 4685, 5120, 5537, 4953, 4536, 4633, 4618, 4569, 4701, 4414, 5345, 6071, 5791, 6110, 6215, 5971, 6110, 5123, 5360, 2484, 0, 512, 0, 1926, 5048, 4729, 5912, 5259, 3980, 4068, 3725, 4185, 5571, 5192, 5748, 7227, 6456, 4796, 3960, 4477, 4503, 5022, 5576, 5856, 6092, 6307, 6193, 6186, 6298, 6258, 6281, 6263, 6282, 6260, 6237, 5530, 4668, 4853, 5218, 5396, 5539, 5622, 5933, 5601, 5723, 5919, 5519, 2740, 63, 89, 0, 152, 0, 473, 0, 3626, 7468, 6547, 6861, 5690, 5245, 4150, 4020, 4716, 4627, 6045, 5836, 8580, 10767, 9753, 6489, 1718, 2213, 1764, 2105, 1754, 2252, 1319, 4565, 8888, 6755, 6164, 5798, 4844, 5279, 5100, 4732, 5260, 4949, 4962, 5070, 4856, 4831, 3854, 3624, 3793, 2801, 710, 0, 132, 0, 268, 0, 2250, 6284, 6344, 6464, 6773, 7657, 7223, 7966, 7181, 8049, 10053, 12092, 21071, 25067, 23972, 24669, 23994, 25035, 20854, 9339, 6839, 8379, 7937, 9113, 9528, 9669, 9030, 9101, 7041, 5569, 5496, 4752, 4778, 4421, 4346, 4256, 4069, 4478, 5150, 5240, 4630, 4825, 3842, 3105, 2594, 1896, 1469, 1212, 465, 576, 2916, 3072, 4205, 5556, 6596, 8035, 8059, 7625, 8116, 7264, 8810, 5747, 15620, 24646, 22339, 22561, 21514, 19532, 19299, 13838, 7544, 10755, 9737, 10510, 8288, 7111, 6446, 4997, 5081, 4491, 4770, 4543, 4140, 4576, 4576, 4237, 3928, 4117, 4558, 4522, 4328, 4289, 2551, 1431, 1957, 1753, 1941, 2477, 3037, 2922, 3115, 3212, 3203, 3189, 3215, 3183, 3228, 3132, 4947, 13790, 14282, 10837, 12989, 12999, 13843, 13418, 12687, 12126, 11121, 10937, 10423, 8714, 8208, 8351, 7329, 6400, 5542, 4618, 4844, 4879, 4622, 4815, 4713, 4705, 4752, 4789, 5589, 5506, 4995, 5218, 4920, 4735, 4570, 4833, 5188, 5113, 5077, 5232, 4903, 5566, 3612, 3459, 5662, 3508, 1995, 1975, 1758, 2386, 3921, 3567, 5369, 5040, 7132, 8687, 4752, 4078, 5290, 6532, 6002, 5458, 5786, 5999, 6371, 6436, 6177, 5601, 4693, 4914, 4588, 4404, 4579, 4838, 4914, 4593, 4424, 4978, 5624, 5295, 5176, 5196, 5186, 5194, 5186, 5199, 5119, 4770, 4742, 5104, 5189, 5443, 5258, 5408, 4302, 2665, 3176, 1486, 3412, 3443, 1225, 1890, 2020, 3760, 4235, 4546, 4887, 3982, 4138, 3839, 2771, 2765, 2515, 2861, 2841, 3689, 4916, 4932, 5542, 5377, 4998, 5085, 4590, 4926, 5239, 5132, 5217, 5115, 5270, 4983, 5883, 6583, 5970, 6213, 6004, 5203, 5102, 5585, 5939, 5499, 5866, 6486, 5757, 5593, 5413, 4085, 1080, 0, 95, 0, 302, 2567, 4936, 3934, 2930, 2917, 3317, 2613, 2317, 3166, 3325, 4273, 4346, 4221, 4329, 4358, 4439, 4767, 5082, 4968, 5058, 4947, 5121, 4796, 5777, 6213, 5254, 5359, 5619, 5936, 6040, 6112, 5843, 5645, 5549, 5842, 6219, 6314, 6631, 6856, 5857, 6725, 6883, 3773, 849, 0, 71, 0, 16, 0, 8, 176, 1799, 2153, 3084, 2162, 3219, 2923, 1387, 3593, 2923, 4356, 5336, 5032, 5246, 5022, 5332, 4791, 6333, 6831, 6052, 6925, 7839, 8972, 8417, 8785, 8276, 7502, 7316, 6708, 6375, 5651, 5993, 6575, 6868, 6596, 6151, 5715, 4879, 3247, 2393, 2377, 2176, 866, 0, 103, 0, 34, 0, 16, 88, 1245, 2164, 1974, 3746, 4765, 4501, 4447, 4816, 3995, 5585, 2357, 13160, 24996, 21107, 19631, 14589, 9649, 5308, 5937, 7208, 8206, 8318, 8175, 8995, 8378, 8325, 6755, 5422, 5172, 4613, 4382, 4796, 5157, 5368, 5269, 5038, 5567, 5148, 5100, 5160, 3631, 2741, 2322, 2354, 1752, 1288, 664, 0, 1521, 2334, 2105, 2255, 2116, 2266, 2046, 2985, 4921, 3446, 15430, 23914, 22600, 23833, 22508, 22093, 20384, 18783, 20385, 13801, 7806, 11603, 10012, 8214, 7829, 8115, 6847, 5678, 5229, 4757, 5353, 5157, 5060, 5056, 5085, 5731, 5544, 5310, 5226, 5211, 4950, 4652, 2843, 1646, 2218, 2157, 2218, 2190, 2195, 2207, 2175, 2326, 2597, 1918, 2097, 2152, 1779, 1814, 1988, 3756, 6440, 8909, 9869, 11077, 11544, 10367, 10541, 10959, 10864, 10646, 10163, 9806, 8748, 8567, 6579, 4810, 5030, 4574, 4743, 4595, 4503, 4746, 4666, 4630, 4587, 5003, 5326, 4845, 5112, 5314, 5282, 5259, 5340, 5170, 5528, 4271, 2564, 2658, 2368, 2363, 2303, 2303, 942, 0, 258, 0, 42, 0, 0, 12, 0, 50, 0, 444, 1286, 2228, 3126, 4292, 4994, 5188, 6564, 6330, 5770, 6010, 5764, 6112, 5538, 6636, 3012, 0, 596, 0, 2026, 4618, 4454, 3908, 4508, 5638, 5966, 4354, 2438, 4382, 1304, 746, 2110, 1460, 2814, 2650, 3090, 3502, 4942, 5782, 5884, 6552, 7054, 7430, 7486, 7462, 8026, 6282, 2572, 0, 5842, 17730, 20206, 21868, 22348, 22206, 22374, 22116, 22548, 21726, 24296, 26202, 24704, 26578, 27254, 25522, 26498, 25866, 24892, 25686, 25530, 26076, 24344, 22824, 25568, 27704, 28442, 29584, 29524, 30178, 30072, 30952, 31708, 30834, 31026, 31088, 30782, 31002, 30854, 30854, 30864, 30170, 29836, 28910, 29690, 25406, 26358, 31060, 29736, 30750, 29652, 31256, 28534, 33834, 16660, 0, 5172, 3860, 7458, 5206, 4240, 4312, 4740, 7612, 4450, 15658, 28284, 26476, 27818, 26742, 26986, 28778, 29956, 29178, 29160, 29702, 30136, 29192, 30148, 27358, 31154, 14878, 22, 5888, 3294, 5270, 4182, 5648, 7822, 5836, 4494, 4642, 4628, 4610, 4700, 4500, 4854, 4604, 11980, 23472, 26864, 27458, 28032, 28960, 29106, 28790, 29320, 30086, 30348, 31422, 32540, 32780, 32926, 33170, 32516, 32830, 32160, 31136, 32080, 31954, 31206, 30864, 29724, 28236, 24720, 25672, 27354, 28312, 18044, 1338, 16106, 30436, 29164, 29554, 29936, 28338, 26114, 26964, 26300, 27100, 25740, 29892, 33530, 31826, 33376, 32734, 31572, 32370, 30236, 33694, 16868, 2502, 6918, 4430, 5528, 4736, 5488, 4998, 6322, 8044, 7990, 8228, 8158, 8148, 8204, 8242, 8112, 7080, 6640, 8390, 6682, 4886, 4552, 3700, 4004, 3922, 3896, 3612, 3798, 3810, 3600, 3736, 3556, 3854, 3286, 5016, 6454, 7504, 8948, 8468, 8866, 8314, 8938, 7346, 6170, 6396, 7558, 8992, 8296, 8094, 8738, 7006, 5160, 5996, 5752, 4920, 4070, 0, 13220, 29662, 25202, 27196, 28294, 28558, 29084, 26208, 25990, 9532, 0, 3592, 0, 708, 0, 190, 0, 120, 0, 352, 0, 2906, 7054, 6108, 6724, 5650, 7134, 8446, 9900, 19734, 26640, 25926, 27340, 25452, 27430, 30050, 27620, 29102, 30862, 27298, 26720, 24600, 28740, 12778, 0, 1584, 0, 398, 0, 0, 294, 0, 2814, 6942, 5866, 6674, 6322, 7686, 9296, 9110, 9258, 9180, 9182, 9286, 9020, 9430, 7474, 9304, 2856, 2420, 4080, 0, 1876, 4982, 8024, 8442, 6830, 7786, 9916, 7510, 7822, 9392, 7784, 6528, 6812, 6932, 7060, 7048, 7334, 6912, 8414, 9682, 9836, 8124, 7256, 6548, 9254, 7044, 17518, 30408, 26020, 26920, 27008, 27216, 27154, 27154, 27166, 27168, 27102, 27414, 28542, 29872, 25522, 26234, 31154, 30766, 32004, 32962, 32772, 31532, 31606, 31624, 31776, 31802, 31166, 31752, 31648, 32420, 31732, 30694, 30108, 29692, 30374, 30680, 31028, 31026, 31050, 31182, 31242, 31446, 31300, 31356, 27672, 24590, 25142, 24994, 26948, 27808, 27868, 27330, 28536, 26206, 30900, 15768, 2846, 9696, 6716, 9382, 9822, 10254, 9026, 7562, 8818, 11638, 24620, 30298, 28252, 28298, 27540, 28782, 28892, 29838, 29706, 30330, 31208, 31828, 32070, 31330, 31760, 28558, 31244, 18110, 5892, 9896, 8370, 9014, 9660, 11014, 10804, 9752, 8700, 9316, 8830, 9492, 8390, 10354, 6478, 19064, 31106, 27320, 30488, 30082, 29922, 29452, 30496, 29594, 29722, 30410, 31016, 31652, 30682, 30922, 31588, 31364, 28514, 29138, 30962, 30048, 30218, 30068, 30694, 31410, 31298, 29548, 30504, 30408, 30844, 31678, 31528, 30674, 29716, 29296, 27026, 29568, 29166, 27466, 28040, 27724, 27938, 27744, 27998, 27574, 28740, 28138, 28742, 29250, 29806, 28790, 30646, 18676, 0, 3916, 8294, 8120, 8504, 9042, 9042, 9852, 10810, 10290, 10574, 10734, 10484, 10418, 10318, 10142, 9550, 10150, 8728, 7674, 7214, 5750, 6790, 5688, 7402, 2074, 2030, 3134, 0, 566, 0, 338, 0, 718, 0, 5588, 12494, 10246, 11260, 10778, 10716, 10938, 9830, 8396, 9710, 10592, 11042, 10150, 10178, 8592, 7272, 8884, 6292, 8168, 2362, 13186, 29444, 27540, 30560, 28780, 28322, 29534, 30082, 28742, 30340, 26914, 29938, 13128, 0, 1632, 0, 464, 0, 124, 0, 158, 0, 554, 0, 4562, 10052, 8480, 9172, 11728, 8794, 19158, 28918, 25434, 27846, 26622, 27890, 28294, 28624, 29130, 28820, 28288, 28082, 27918, 25474, 28158, 24454, 28880, 13622, 0, 1680, 0, 248, 192, 0, 3706, 9138, 8528, 9306, 9334, 8894, 10334, 11798, 11196, 11380, 11496, 11008, 12062, 10094, 13776, 3128, 9382, 31212, 10342, 0, 1602, 0, 4892, 5496, 0, 6426, 12040, 9460, 10538, 10608, 10962, 10186, 10094, 11024, 10602, 10508, 10918, 10614, 11606, 12156, 12316, 11120, 10452, 8982, 12548, 9322, 19418, 30172, 26450, 29688, 28036, 28786, 28946, 28944, 28904, 29036, 28722, 29360, 27776, 28974, 28500, 27834, 30960, 30184, 31744, 33186, 32462, 31816, 32034, 32232, 32346, 31908, 31438, 31678, 31992, 31640, 31960, 30782, 29280, 29602, 29942, 30246, 31150, 30240, 30550, 30998, 30286, 30366, 30164, 30782, 29272, 28310, 27212, 25630, 26130, 26926, 26860, 27116, 26608, 27558, 25810, 29290, 17954, 6940, 10570, 9182, 11936, 12068, 12472, 10504, 9910, 9418, 12224, 10106, 17534, 31026, 28490, 28698, 29390, 29844, 30346, 30488, 31116, 31400, 32364, 32320, 31706, 32806, 30716, 32256, 18774, 8150, 12196, 10690, 11516, 11012, 11294, 11160, 10532, 10744, 11514, 11050, 11670, 10638, 12474, 8858, 20598, 31838, 28196, 30672, 30244, 30044, 29686, 28972, 29502, 30422, 29974, 30878, 31582, 29590, 29116, 30454, 30832, 31958, 27804, 28882, 32478, 29236, 29762, 30562, 28988, 29918, 29540, 30640, 30310, 29534, 30608, 30134, 31452, 30210, 29212, 29846, 29346, 29342, 29378, 29376, 29366, 29408, 29302, 29516, 29140, 30352, 29172, 29110, 28880, 25572, 27914, 28300, 29766, 17970, 8590, 11170, 9832, 10626, 10548, 10682, 11894, 12510, 12146, 10714, 9106, 9640, 9706, 10752, 12178, 9546, 7856, 9082, 9584, 9840, 9280, 8234, 6726, 8468, 3472, 0, 412, 0, 156, 0, 206, 0, 638, 0, 5140, 11786, 10966, 12996, 12308, 12250, 12816, 11576, 10612, 10310, 11072, 11430, 9690, 8920, 10132, 10620, 10980, 9928, 10840, 6960, 16180, 29194, 27482, 29498, 28984, 29276, 29416, 29372, 29080, 29476, 25898, 28774, 12012, 0, 1456, 0, 400, 0, 0, 140, 0, 650, 0, 5214, 11206, 9802, 9698, 14532, 19218, 24944, 28570, 26836, 29310, 29186, 29682, 29106, 28988, 29752, 30922, 30824, 31118, 30492, 29216, 28804, 29344, 27696, 29128, 24476, 32678, 9974, 8764, 14326, 0, 2996, 0, 5612, 11434, 10380, 11542, 10908, 12046, 12788, 12556, 12652, 12652, 12524, 12872, 12092, 13184, 9740, 15238, 23358, 28644, 12396, 0, 1710, 0, 1104, 0, 5548, 12374, 10256, 11400, 11170, 11372, 10802, 11208, 11522, 11436, 11790, 12096, 11664, 12322, 13444, 13006, 12076, 12328, 11470, 12898, 9190, 20246, 29512, 27104, 31168, 30394, 31554, 31524, 31472, 31704, 31234, 32140, 29276, 27630, 31270, 28394, 27214, 30204, 29960, 31636, 33238, 32478, 32002, 32230, 32682, 32376, 31678, 31042, 31848, 32110, 31510, 30926, 30232, 29994, 30256, 30686, 31222, 31036, 30614, 29934, 29528, 29408, 30386, 30776, 29480, 25718, 26286, 25280, 24012, 26088, 25844, 27132, 25942, 27742, 24624, 30664, 12098, 1146, 12038, 8726, 11878, 11898, 12368, 10326, 11072, 10178, 12236, 9404, 19874, 32322, 28184, 29194, 30020, 30982, 30824, 30626, 29804, 30562, 31808, 31832, 32010, 31140, 31398, 28808, 30458, 18444, 8748, 12384, 10476, 11890, 11690, 11442, 11312, 11966, 12530, 12180, 12690, 11808, 13398, 10244, 20584, 31274, 29166, 31202, 30238, 31220, 31422, 31504, 31858, 31040, 32182, 29786, 30518, 30430, 27714, 29872, 28022, 28068, 26102, 24290, 28730, 30826, 29872, 30316, 31400, 31746, 32026, 32858, 33006, 31474, 29698, 30174, 30682, 30156, 30762, 30982, 30364, 29814, 29478, 29590, 29522, 29572, 29528, 29600, 29138, 27788, 29262, 27468, 24176, 26748, 24974, 28774, 28256, 31556, 12454, 0, 2440, 3768, 13398, 10038, 12688, 12962, 12806, 11492, 10478, 10476, 11168, 12468, 11526, 9194, 9736, 11000, 11286, 11002, 9430, 11080, 7788, 15668, 32418, 14914, 0, 14988, 29556, 25866, 27326, 27112, 26136, 28944, 18952, 9072, 11918, 11594, 13356, 12628, 11714, 10650, 11168, 10196, 12048, 10820, 7808, 8744, 9772, 10904, 10108, 10720, 7668, 16266, 30326, 31432, 31752, 30982, 31698, 33292, 32516, 33860, 32082, 30946, 26702, 30178, 13420, 0, 1674, 0, 474, 0, 130, 0, 252, 0, 1106, 0, 6816, 7354, 19052, 9162, 8886, 30754, 25134, 30210, 29000, 30636, 30522, 30378, 30106, 31992, 31742, 31816, 31734, 31168, 29062, 27994, 28356, 28222, 24542, 31124, 10350, 7412, 32202, 9330, 0, 0, 3922, 10920, 9308, 11190, 10730, 10342, 11998, 12826, 12318, 12606, 12270, 12842, 11782, 13826, 9106, 17330, 25862, 30038, 13926, 0, 1634, 0, 0, 794, 0, 6578, 6360, 48, 11722, 2844, 4016, 11864, 9820, 11236, 10160, 11074, 11118, 11332, 11246, 12378, 12524, 10652, 12272, 8668, 17568, 27964, 27404, 29372, 30088, 31050, 30686, 31224, 31140, 31216, 31130, 31250, 31044, 31472, 29766, 26406, 27014, 29542, 29706, 31584, 33282, 32756, 33008, 32632, 33020, 33272, 32464, 32048, 32052, 32322, 32694, 31174, 30182, 30086, 31154, 31186, 30922, 32054, 32264, 32446, 31256, 29596, 30544, 31742, 29058, 29380, 27150, 24752, 26288, 25462, 25730, 26658, 27052, 27160, 26732, 27624, 25938, 29326, 18200, 7222, 11620, 10304, 11994, 10180, 11650, 8212, 19794, 30978, 27128, 29258, 29408, 30726, 31052, 31604, 31126, 30642, 31204, 33446, 33594, 33114, 32424, 32930, 32868, 33462, 30462, 31786, 19136, 7508, 12684, 10992, 11842, 11518, 11870, 11688, 11496, 11418, 11318, 11134, 11634, 10632, 12512, 8740, 21192, 33918, 29718, 31660, 30758, 30190, 32376, 32178, 32820, 33720, 27874, 29558, 33428, 29386, 30350, 32562, 28756, 25258, 23718, 28050, 30882, 30386, 30188, 30644, 31646, 30840, 31494, 31930, 31830, 30832, 30130, 30028, 30500, 31512, 31014, 30708, 30948, 30256, 29538, 29772, 29616, 29786, 29522, 29994, 28980, 30122, 26702, 24152, 24656, 26718, 26838, 28716, 15084, 0, 4046, 8366, 10170, 10720, 11404, 10898, 12198, 11992, 10556, 10562, 9864, 9670, 9348, 8830, 7896, 8182, 8726, 9476, 9776, 8378, 6760, 8786, 3852, 0, 470, 0, 136, 0, 68, 0, 202, 0, 708, 0, 5584, 11954, 9420, 10998, 10162, 10192, 11000, 11672, 10834, 9788, 9912, 9612, 8774, 9724, 8914, 9910, 7586, 11252, 724, 12692, 33166, 28230, 31110, 30242, 32048, 33430, 30470, 30350, 32412, 30112, 28416, 28940, 21060, 4156, 0, 260, 0, 62, 0, 0, 104, 0, 458, 0, 4278, 10958, 5540, 0, 11382, 26552, 25444, 28816, 28116, 29338, 28612, 28200, 29142, 31754, 30242, 27528, 30494, 29866, 29710, 28396, 27446, 28152, 25248, 30916, 12758, 0, 1678, 0, 990, 0, 4450, 9522, 8420, 9806, 10134, 10168, 10762, 11900, 11366, 11714, 11320, 11950, 10842, 12908, 8044, 16716, 29484, 22016, 6710, 0, 586, 0, 0, 836, 0, 6140, 6048, 0, 626, 56, 0, 4470, 10954, 9716, 10700, 10034, 10496, 10446, 10686, 10772, 11258, 10760, 11930, 8900, 16892, 27360, 27440, 30392, 29082, 29900, 30916, 30650, 30894, 30780, 30818, 30826, 30772, 30940, 29826, 25772, 26884, 31168, 30556, 32364, 34144, 33314, 33726, 33354, 33350, 32510, 31616, 31424, 31418, 31820, 31224, 31444, 30552, 30250, 31224, 30474, 30498, 31364, 31782, 31578, 30736, 29752, 31090, 28016, 25206, 27040, 27336, 26326, 25328, 26480, 27946, 30682, 32432, 31352, 32886, 30280, 35334, 19042, 3852, 10556, 9056, 10714, 9426, 9622, 9654, 8960, 9202, 10548, 21094, 28462, 27992, 29644, 29348, 29794, 30404, 31546, 31792, 32676, 33096, 32570, 32428, 31010, 32578, 29180, 31760, 14238, 0, 6386, 10096, 9512, 10154, 10362, 10246, 10018, 9536, 9744, 9464, 10032, 8968, 10926, 7022, 19842, 32844, 29122, 31852, 30314, 31326, 31226, 31856, 31252, 32272, 30378, 27150, 29356, 28890, 28816, 29752, 27346, 24882, 24592, 28664, 31080, 29762, 30032, 29650, 30324, 30398, 31246, 30532, 29496, 29258, 28532, 28746, 29022, 29600, 30118, 30268, 30006, 29734, 29668, 29576, 29604, 29594, 29592, 29616, 29370, 27844, 26178, 25046, 27324, 29388, 31072, 26350, 29650, 13440, 0, 2138, 0, 4420, 9644, 9328, 9048, 8416, 9024, 8682, 8722, 8902, 8712, 8596, 7362, 7482, 8544, 8718, 8194, 8172, 3228, 0, 1014, 0, 2434, 0, 15306, 15258, 0, 2246, 0, 344, 256, 0, 4564, 10384, 8438, 9146, 9008, 9436, 8906, 8960, 8608, 8998, 7352, 5708, 6842, 6794, 8672, 6874, 9590, 0, 11996, 31096, 28736, 31354, 30560, 31456, 31462, 30604, 30698, 30180, 30106, 27354, 30994, 13704, 0, 2004, 0, 1576, 0, 8938, 19884, 16616, 18130, 17574, 17356, 18584, 13476, 3730, 0, 8450, 24366, 26326, 28426, 28624, 29746, 29362, 28042, 29814, 32492, 32020, 31390, 32174, 30036, 30218, 28060, 27790, 29040, 28184, 27500, 26188, 9120, 0, 874, 0, 0, 1874, 4952, 5902, 7106, 7440, 8394, 7904, 8726, 8262, 7600, 7666, 7934, 7206, 8730, 5572, 15348, 23764, 28798, 13538, 0, 1736, 0, 486, 0, 88, 0, 0, 48, 0, 164, 0, 1672, 5718, 6848, 7396, 7524, 7756, 8416, 8946, 8554, 9278, 7630, 10976, 978, 10330, 27202, 24462, 28128, 27834, 28864, 29102, 29972, 30482, 31088, 30950, 30908, 31116, 30672, 31608, 28202, 23846, 28852, 31832, 32656, 33806, 33120, 33260, 32804, 32842, 33792, 33806, 32472, 32342, 32468, 32384, 32138, 31790, 31018, 31550, 31752, 30700, 31700, 31536, 31846, 31502, 30894, 30308, 28054, 25796, 28380, 30164, 26644, 26420, 26816, 31418, 32252, 29998, 31062, 30904, 30320, 31878, 28764, 35072, 14810, 0, 7376, 5298, 6864, 6326, 5304, 10820, 22934, 26930, 27964, 28882, 29340, 29590, 29540, 29804, 30938, 30312, 31644, 32076, 32510, 32616, 30796, 32078, 28844, 31416, 13386, 0, 4024, 5796, 7600, 7878, 8232, 8016, 8086, 7564, 6306, 6136, 6500, 6138, 6762, 5630, 7694, 3582, 17196, 31776, 28216, 30978, 30772, 31660, 31944, 32330, 30184, 28064, 28024, 27846, 31028, 28974, 25974, 27430, 26156, 31124, 32712, 30180, 31582, 31564, 31668, 31278, 31426, 32140, 30832, 30048, 29944, 28720, 28958, 29458, 29802, 29250, 30890, 31724, 32726, 29832, 26286, 27358, 26910, 26992, 27228, 26566, 28746, 28746, 289, 0, 4256, 4826, 10812, 17042, 14653, 15511, 15111, 15826, 15465, 15130, 14698, 15256, 14737, 17222, 10234, 4451, 6847, 7899, 8902, 7273, 7890, 7604, 7693, 7783, 7449, 8401, 7821, 8501, 4392, 13281, 14206, 6084, 9766, 7507, 7631, 7117, 6911, 7133, 8017, 7990, 7919, 8004, 7173, 6954, 5216, 4964, 2271, 0, 310, 0, 170, 0, 321, 0, 2852, 8105, 8511, 13690, 19412, 10621, 4878, 5193, 4573, 6474, 5667, 6187, 5723, 6316, 5264, 8760, 12912, 11409, 11704, 11666, 10363, 10113, 12146, 13504, 13358, 13510, 12826, 10840, 8462, 7106, 4284, 2921, 3586, 3527, 4203, 4355, 4501, 4111, 3992, 3646, 4542, 4863, 3164, 912, 0, 118, 0, 142, 0, 412, 0, 3438, 8845, 8051, 8871, 7930, 9332, 6710, 15525, 27258, 27619, 28549, 28158, 30449, 27965, 25281, 22522, 23790, 17926, 13264, 14150, 12732, 15037, 13784, 14901, 14825, 14333, 13377, 12535, 11680, 9519, 6927, 4537, 4653, 3476, 1777, 519, 331, 172, 2206, 2878, 1804, 3033, 5972, 4255, 1383, 2774, 2239, 2786, 2066, 3234, 1022, 7636, 10582, 5607, 7477, 7419, 9558, 7557, 18013, 27002, 25056, 25745, 24128, 23948, 24807, 23501, 23153, 23239, 26964, 20142, 13520, 17526, 14629, 14662, 13754, 12493, 12404, 10920, 8079, 8210, 8140, 6619, 6976, 6434, 6130, 5205, 3934, 2952, 3117, 3459, 3172, 3408, 3084, 3625, 2577, 5989, 9467, 8927, 9627, 10369, 9381, 7444, 7558, 7235, 8419, 7337, 12067, 18005, 18869, 19401, 17937, 18593, 19135, 20043, 18615, 13822, 16225, 17397, 15313, 15568, 16068, 17344, 16797, 15216, 10708, 7401, 6859, 7004, 6441, 5476, 6151, 6270, 5525, 5246, 5321, 5258, 5341, 5206, 5471, 4470, 2426, 2005, 2668, 5485, 7245, 7357, 7948, 7790, 7972, 8175, 8330, 9090, 9612, 10064, 10358, 7972, 7729, 11607, 15294, 17134, 14927, 12849, 10880, 9609, 10037, 10295, 12146, 12324, 12289, 10351, 7805, 8809, 10439, 12640, 8895, 5556, 5517, 4600, 4953, 4800, 4824, 4913, 4666, 5496, 6295, 6525, 6628, 5252, 5731, 6151, 5180, 5701, 6679, 6799, 7063, 6835, 5865, 5864, 7408, 8253, 8662, 9323, 9552, 7858, 7575, 6555, 12090, 17765, 15333, 17607, 11520, 5849, 9343, 11495, 6154, 1460, 2498, 2110, 1112, 393, 1026, 1066, 1020, 1168, 867, 1434, 294, 4093, 8022, 5821, 5415, 5333, 5594, 6258, 6794, 6544, 6216, 5829, 5917, 6705, 7373, 6569, 7119, 7886, 6732, 6600, 6621, 6690, 7596, 7752, 8609, 9187, 8277, 7742, 6003, 2017, 0, 0, 81, 284, 5601, 8166, 13505, 10478, 3504, 5690, 4572, 5153, 4885, 4947, 5049, 4579, 4139, 3721, 3929, 4581, 4892, 7108, 7409, 10041, 12381, 12964, 11878, 9780, 10536, 8073, 6311, 6469, 6538, 7012, 6280, 6430, 3191, 827, 2294, 2004, 3888, 4183, 4719, 3877, 7257, 8456, 3790, 1326, 0, 169, 0, 39, 0, 35, 0, 156, 0, 560, 0, 4260, 8421, 7034, 6713, 5820, 6916, 8369, 10451, 14137, 8322, 5696, 11862, 11815, 13687, 12752, 10777, 9671, 10350, 11744, 12296, 13189, 10919, 10127, 10459, 9901, 9051, 7451, 6115, 4695, 5105, 4680, 4885, 5383, 3973, 2671, 2144, 3146, 3127, 2121, 2498, 2259, 2467, 2215, 2645, 1208, 34, 4545, 8037, 7819, 7321, 7749, 8231, 6092, 8616, 15556, 22752, 27753, 27748, 27355, 25871, 24054, 21311, 14076, 14767, 14511, 11611, 13717, 13681, 13537, 14217, 15397, 14662, 14449, 12499, 10846, 8997, 6944, 6258, 5024, 4517, 4460, 2728, 1656, 1876, 1919, 1619, 2293, 916, 4746, 3509, 0, 325, 63, 0, 3040, 8845, 8353, 10638, 10695, 7906, 8044, 8017, 9105, 8713, 14642, 24441, 25049, 22816, 20539, 18879, 16797, 14384, 12138, 11859, 12473, 13311, 15043, 14706, 14804, 13085, 10783, 10492, 9541, 8590, 9273, 8195, 6817, 7262, 7005, 7208, 6980, 7346, 6266, 4849, 2778, 2773, 5677, 6529, 7166, 7732, 8467, 8198, 8795, 9425, 8862, 8000, 7566, 7217, 8127, 9639, 9797, 10441, 13031, 17775, 18706, 19598, 15524, 15861, 17478, 14166, 14548, 13789, 14896, 15305, 15091, 14720, 14047, 15126, 15300, 12208, 10964, 11300, 11040, 11363, 10861, 11805, 8693, 5234, 6981, 7497, 8167, 6911, 6042, 6414, 5745, 5256, 5674, 6442, 7019, 7167, 6992, 7787, 8342, 8481, 9068, 8652, 9161, 9501, 9239, 8516, 7400, 8706, 9874, 10950, 11837, 12006, 9749, 14706, 13483, 8689, 10536, 9213, 8936, 8182, 8290, 8245, 8230, 8293, 8169, 8431, 7421, 5401, 4867, 5008, 4978, 5064, 5554, 5844, 6121, 6206, 6392, 6590, 6281, 6674, 7180, 6189, 5778, 6392, 6652, 6444, 6633, 6304, 6819, 7971, 6789, 7220, 7555, 9029, 10196, 8475, 8141, 8978, 10116, 9486, 8935, 8927, 8266, 8086, 8110, 8144, 8042, 8255, 7844, 8674, 6027, 3821, 4357, 4494, 4522, 4695, 6461, 7760, 8384, 7947, 7188, 6209, 5659, 6041, 7089, 6794, 6993, 6512, 7298, 7186, 7654, 9190, 7810, 7490, 7554, 7580, 7671, 7226, 7913, 8402, 8172, 8582, 8459, 8439, 7599, 7452, 5125, 781, 0, 0, 125, 0, 498, 0, 3767, 6901, 4966, 5439, 4097, 4735, 4984, 6161, 6826, 6449, 5791, 5250, 5592, 6318, 6032, 6829, 7260, 7870, 8941, 9267, 9085, 8710, 8632, 8185, 7225, 6921, 7507, 7012, 6556, 6750, 6519, 6399, 7067, 7610, 7437, 7797, 7673, 7041, 7048, 7090, 6927, 7273, 6612, 7939, 3552, 0, 560, 0, 1390, 4822, 8296, 9033, 8774, 8434, 6062, 6037, 5386, 4626, 6186, 6598, 6680, 7577, 6040, 4401, 8026, 10260, 9808, 11101, 9915, 8347, 9973, 11020, 11003, 11521, 12496, 10336, 8956, 8750, 7217, 7012, 6317, 6135, 6242, 6209, 6205, 6256, 6136, 6389, 5611, 4713, 2592, 149, 16, 8, 0, 144, 0, 1437, 4689, 7038, 7886, 8636, 8943, 8747, 7509, 9955, 12482, 14843, 23422, 27284, 26873, 25422, 25275, 24647, 24883, 18095, 17252, 14630, 9853, 13175, 12309, 12614, 12481, 14053, 14432, 13410, 13068, 12956, 13324, 12574, 14109, 9137, 4683, 5988, 5518, 6164, 5714, 6219, 6000, 5499, 5280, 5821, 6981, 4091, 607, 0, 1961, 6452, 8050, 9351, 9461, 9672, 9089, 8369, 8695, 8961, 9616, 12255, 17000, 21080, 22186, 21433, 21174, 18024, 16143, 13759, 10828, 11751, 12252, 13377, 14009, 13705, 14077, 13492, 14601, 10940, 6676, 7426, 6335, 5782, 5314, 5344, 5592, 5377, 5152, 5423, 5603, 5248, 4482, 1868, 3000, 6673, 8334, 9184, 9251, 8841, 8109, 8453, 8422, 8749, 9036, 9271, 10083, 10532, 10908, 11122, 13071, 18361, 22297, 18131, 15557, 15652, 15794, 16557, 15772, 16037, 16003, 15830, 16314, 14564, 12049, 10361, 8334, 7504, 6755, 6151, 5654, 5733, 5829, 6033, 6054, 5570, 6788, 7736, 7750, 6673, 5591, 5899, 5329, 5559, 5591, 5640, 6377, 6077, 7172, 8901, 9427, 10062, 9867, 9676, 9431, 9193, 9406, 8601, 10682, 11086, 15234, 19352, 18149, 18624, 18601, 18188, 19275, 15558, 12716, 15368, 13002, 10310, 9572, 8344, 7682, 8076, 7481, 6042, 5405, 5125, 5179, 5242, 5063, 5402, 5229, 5825, 6035, 6172, 6648, 6707, 8108, 7880, 5941, 5972, 6432, 6940, 5908, 5110, 4514, 5560, 7152, 6465, 6614, 6819, 8894, 10231, 9862, 10030, 9967, 9946, 10082, 9436, 8112, 8764, 10022, 8326, 5514, 6301, 5451, 4049, 3873, 3515, 4266, 4641, 4217, 4877, 6657, 6916, 6985, 7146, 6293, 5285, 5292, 4708, 4975, 5312, 5188, 5129, 6127, 7046, 6456, 6824, 6987, 6407, 6434, 6806, 6920, 7112, 7589, 7803, 7763, 7763, 7783, 7740, 7857, 6849, 1734, 0, 0, 1971, 4751, 9430, 11265, 8010, 6308, 4572, 4962, 4702, 5209, 4797, 4975, 5197, 5384, 5280, 4772, 4821, 5135, 5160, 5626, 6681, 6890, 6944, 7206, 7505, 8015, 8218, 8009, 8442, 7666, 7899, 7999, 7234, 6507, 5554, 5853, 5737, 5744, 5836, 5604, 6387, 7157, 7200, 8151, 3767, 0, 164, 0, 21, 24, 0, 186, 0, 1977, 6951, 8538, 8066, 7582, 7017, 6644, 5193, 4000, 5631, 5835, 7245, 6450, 4315, 4840, 6801, 9319, 9842, 9803, 7954, 7790, 8675, 9140, 9835, 9499, 9425, 9481, 9351, 9610, 9129, 10076, 7140, 5341, 7151, 6285, 6160, 5458, 5524, 6156, 5978, 5471, 3383, 513, 0, 0, 52, 0, 212, 0, 2155, 7065, 7698, 8623, 8669, 9508, 10534, 8965, 8525, 8566, 17632, 25044, 23188, 23363, 22768, 22618, 20107, 16400, 16916, 12124, 8459, 9475, 9054, 9129, 9374, 8679, 10851, 10312, 5593, 6312, 6670, 5840, 5434, 5269, 4962, 4860, 5042, 5277, 5128, 4632, 3425, 3277, 3485, 5696, 7826, 4451, 0, 2051, 5446, 7110, 8543, 8812, 10306, 11035, 11441, 9740, 9913, 9422, 11962, 11357, 16812, 23041, 21910, 22839, 21354, 22062, 21520, 22145, 21173, 23020, 17085, 11305, 12181, 10771, 10632, 8359, 8131, 7334, 6743, 7715, 6642, 5734, 6019, 6187, 6143, 5312, 4902, 5387, 4339, 4417, 4078, 2948, 1685, 3883, 7619, 7767, 8484, 8423, 8234, 7997, 7926, 8449, 8614, 9975, 11611, 11250, 11964, 12911, 12958, 12955, 13009, 12875, 13140, 12609, 14261, 15150, 13526, 13650, 12801, 11874, 10339, 9958, 8384, 6692, 7000, 6379, 6339, 6674, 5930, 6036, 6250, 5103, 4484, 5245, 6337, 5814, 4644, 4131, 4288, 3652, 3444, 3382, 3596, 3991, 4950, 3140, 5165, 8340, 7939, 8500, 8285, 8736, 8631, 8648, 8718, 8538, 8897, 8161, 10523, 12560, 12316, 12263, 13535, 11760, 8523, 10261, 11176, 10292, 8730, 9119, 7424, 6372, 7126, 7131, 6535, 5618, 5964, 5240, 4419, 4742, 4497, 4551, 4924, 4996, 5137, 4781, 4606, 4753, 4455, 4276, 4554, 4791, 5499, 5462, 4925, 4844, 4694, 4750, 4722, 4741, 4716, 4758, 4796, 6182, 7536, 8737, 6268, 5957, 8596, 6950, 7500, 5725, 5131, 5581, 4918, 5467, 4827, 3872, 3493, 4081, 4088, 4045, 4621, 5923, 6208, 7116, 6465, 5803, 5505, 5298, 5412, 5086, 5284, 5307, 5097, 5115, 5638, 5365, 5510, 5797, 5852, 5840, 5858, 5823, 5890, 5755, 6192, 6618, 6604, 6400, 5902, 5730, 4878, 3551, 1887, 471, 0, 1003, 3844, 4726, 5212, 5564, 4915, 4658, 4298, 3889, 4234, 4436, 5294, 5712, 5710, 5019, 4107, 4654, 4556, 4487, 5211, 5859, 5744, 6611, 7776, 8546, 6960, 5759, 6280, 6051, 6164, 6119, 6111, 6179, 5881, 5371, 5384, 5517, 5558, 5897, 6538, 5589, 7718, 7422, 10029, 0, 22043, 20249, 0, 2987, 0, 624, 18, 0, 3514, 8723, 8553, 8778, 6121, 4815, 4425, 4269, 4312, 4999, 6362, 5429, 3201, 2255, 2581, 2375, 3625, 6078, 6375, 6363, 6401, 6304, 6498, 6112, 7291, 7781, 6165, 5222, 4619, 4952, 4630, 4641, 5061, 5276, 5239, 5424, 5388, 4046, 3067, 3665, 2681, 1797, 847, 0, 69, 22, 0, 285, 0, 2570, 6612, 6377, 6927, 7155, 8070, 8995, 9462, 9186, 8151, 15052, 23555, 24252, 24062, 24262, 23811, 24693, 23056, 26305, 15754, 5766, 9943, 8286, 10119, 9728, 11510, 10363, 7652, 6742, 4655, 4841, 4344, 3762, 3847, 3890, 3717, 4022, 5031, 4536, 5096, 3629, 2314, 2794, 1932, 2009, 1717, 1138, 671, 2973, 5319, 4745, 6516, 7210, 8481, 11041, 9274, 9346, 9939, 9982, 9582, 10471, 8574, 15343, 23780, 17280, 13866, 11384, 9381, 11536, 10656, 10736, 10898, 11206, 9125, 6751, 6610, 5270, 5197, 4571, 4594, 4705, 4519, 4443, 4594, 4631, 4356, 4088, 4103, 4044, 4203, 2680, 1505, 1971, 1907, 2125, 1839, 3319, 5651, 5351, 6783, 7340, 6491, 6812, 6636, 6754, 6637, 6849, 8004, 13639, 14672, 13325, 14761, 15756, 16061, 15357, 13901, 12315, 13128, 11341, 9186, 8141, 7610, 7129, 6523, 6792, 5852, 4956, 4881, 4492, 4872, 5206, 5495, 4694, 4414, 4997, 4640, 4802, 5123, 4840, 4296, 4173, 4097, 4612, 5493, 4913, 4349, 4533, 4413, 4524, 4358, 5088, 6723, 3804, 1411, 1805, 1681, 1559, 2033, 1901, 3459, 5025, 5090, 7006, 4974, 3547, 5018, 5405, 5468, 5246, 5489, 5882, 6323, 6431, 6451, 5372, 4553, 4641, 4660, 4917, 4470, 4385, 4411, 4724, 4640, 4452, 4431, 4457, 4491, 4401, 4430, 4426, 4407, 4455, 4358, 4651, 4896, 5284, 5794, 5013, 4768, 4062, 2724, 2160, 1797, 1454, 1165, 1276, 1143, 1281, 994, 2047, 3590, 3447, 3026, 3816, 4019, 2696, 2572, 2826, 3075, 2979, 3528, 4134, 4830, 5590, 5649, 5465, 5120, 5244, 5124, 5256, 5711, 5815, 5801, 5804, 5806, 5798, 5815, 5797, 5993, 5924, 5709, 5666, 5546, 5957, 5479, 5807, 6433, 5917, 5439, 5107, 4765, 3838, 2040, 244, 88, 635, 917, 2858, 4050, 3012, 1407, 1929, 3649, 2551, 2099, 2792, 3510, 4454, 4919, 4775, 4496, 4131, 4074, 4498, 4996, 5190, 5137, 5170, 5137, 5185, 5101, 5310, 5147, 4885, 4937, 5209, 5546, 5348, 5011, 4957, 4937, 4899, 5537, 5714, 5799, 5777, 6087, 5270, 4747, 2002, 0, 208, 0, 59, 0, 6, 1, 101, 1486, 2924, 4760, 2121, 3026, 2289, 2889, 4493, 2477, 5354, 5225, 5212, 5163, 5219, 5123, 5310, 4915, 6350, 8530, 8399, 9082, 8716, 7956, 6363, 5250, 4780, 4055, 4232, 3872, 4139, 3885, 3701, 3891, 4092, 4118, 3897, 3373, 2814, 2709, 2241, 2466, 1790, 247, 0, 0, 8, 0, 44, 0, 395, 1097, 1624, 1405, 2197, 5170, 6221, 5807, 6353, 5444, 7045, 3915, 14138, 23608, 16167, 16561, 9979, 3967, 5995, 7213, 8494, 9075, 9365, 9796, 8907, 8329, 7137, 5526, 5846, 5580, 4705, 4300, 4553, 4698, 4004, 3569, 3816, 3831, 3634, 3741, 2047, 871, 1309, 1095, 1233, 482, 0, 18, 403, 1123, 1160, 1142, 1228, 1021, 1438, 616, 2842, 3890, 11564, 21085, 22558, 21513, 21237, 17594, 18296, 10432, 3685, 9136, 8068, 10724, 9848, 8577, 7705, 6582, 6394, 5979, 5378, 5234, 5587, 5535, 5082, 5465, 5812, 5496, 4832, 4382, 4635, 4982, 4597, 4398, 2931, 1727, 2155, 2138, 2258, 2182, 2275, 2111, 2421, 1824, 3253, 2030, 2852, 3328, 1416, 3887, 3510, 5172, 7602, 6866, 9957, 12655, 12566, 12222, 11215, 9535, 9115, 9935, 9238, 9525, 8018, 7228, 6238, 5014, 5062, 5077, 5143, 4922, 4597, 4460, 4362, 4080, 4188, 4450, 4256, 4491, 5090, 5035, 5080, 5058, 5065, 5066, 5058, 5090, 5090, 12459, 12423, 12535, 12532, 12763, 12474, 12599, 13049, 13006, 12654, 12724, 12635, 11908, 12638, 11716, 12948, 5370, 0, 811, 0, 1026, 0, 3033, 0, 19765, 19920, 0, 4649, 1500, 0, 14921, 34292, 8741, 0, 652, 0, 235, 0, 96, 0, 123, 0, 442, 0, 3635, 8725, 9523, 10761, 11382, 10918, 12667, 5334, 0, 0, 3353, 10998, 11377, 11564, 12322, 12704, 12303, 13039, 12944, 13161, 12780, 13467, 12211, 14713, 6510, 0, 828, 0, 329, 0, 392, 0, 2750, 6176, 5540, 6035, 5570, 5525, 4278, 1277, 0, 114, 0, 0, 77, 0, 335, 0, 3373, 11215, 13016, 13917, 14293, 14715, 14953, 15152, 15578, 15639, 15587, 14784, 14377, 14565, 14632, 14641, 14607, 14671, 14564, 14760, 14104, 13345, 12411, 3861, 0, 394, 0, 115, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 32, 0, 158, 0, 552, 0, 5036, 14847, 16341, 16862, 15945, 16129, 16391, 16281, 16398, 16573, 16537, 16497, 16652, 16301, 16992, 15611, 17445, 7114, 0, 414, 364, 0, 6938, 17219, 15414, 15870, 15787, 13525, 13543, 5825, 0, 701, 0, 106, 73, 0, 617, 0, 5248, 12794, 12756, 15220, 15055, 15384, 15543, 16040, 16677, 17094, 17213, 17373, 17459, 17387, 17188, 17077, 17111, 17086, 17114, 17072, 17151, 16932, 16676, 16793, 16413, 17194, 15904, 17946, 6928, 0, 0, 4855, 15577, 15785, 16737, 16852, 17047, 17035, 17198, 17132, 17241, 16272, 15052, 15100, 14675, 14658, 14986, 14765, 14810, 14921, 14829, 14472, 14442, 14379, 14126, 10692, 11940, 14746, 13992, 14570, 14259, 14472, 14271, 14547, 14042, 15656, 17156, 16540, 16339, 16217, 16436, 16217, 16500, 16594, 16196, 15131, 14804, 14670, 14539, 15675, 16380, 16736, 16710, 16803, 16696, 16337, 16391, 16633, 16899, 16757, 17225, 17247, 17424, 16949, 16496, 16076, 14227, 14079, 13535, 13105, 13250, 13392, 13568, 13527, 13125, 14062, 12259, 15790, 5411, 3809, 15233, 6397, 9943, 14900, 13722, 14631, 14547, 14947, 14825, 14917, 14899, 14503, 15087, 14223, 15894, 7850, 0, 7627, 15279, 14274, 15825, 15509, 15846, 15939, 16257, 16319, 16273, 16322, 16528, 16474, 16431, 16262, 15898, 16050, 11934, 7549, 6769, 6313, 6524, 6370, 6518, 6306, 7283, 10421, 10742, 14402, 6411, 0, 796, 0, 230, 0, 47, 0, 0, 19, 0, 88, 0, 302, 0, 3355, 12744, 15820, 15930, 16227, 16321, 16510, 17113, 16997, 16649, 15282, 15013, 15878, 16170, 16750, 16536, 16896, 17344, 17513, 17001, 16883, 16633, 17216, 16085, 18377, 10740, 2480, 4209, 3642, 3857, 3779, 4028, 10579, 5568, 0, 0, 1629, 0, 19222, 17035, 0, 4099, 0, 4274, 0, 19338, 26646, 148, 1159, 0, 378, 0, 184, 0, 504, 0, 4511, 12413, 14706, 17255, 17345, 17954, 18100, 17684, 17194, 17331, 17275, 17282, 17329, 17104, 16870, 17106, 17003, 16512, 17030, 14486, 9682, 9441, 9623, 10216, 9126, 11650, 5533, 0, 572, 0, 0, 942, 367, 25059, 17884, 0, 5866, 0, 17843, 26282, 2516, 303, 0, 23, 171, 0, 741, 0, 6307, 17050, 17252, 18277, 17774, 18079, 17843, 18116, 17645, 19132, 20442, 19636, 20074, 18737, 17330, 18183, 18792, 19282, 20272, 20599, 20422, 20400, 19657, 19866, 17318, 19309, 8112, 0, 666, 67, 0, 5438, 14993, 11098, 11972, 13467, 4160, 0, 402, 0, 120, 0, 28, 0, 0, 0, 0, 77, 0, 385, 0, 1347, 0, 10800, 24232, 20184, 22444, 20767, 20897, 20321, 20368, 20617, 20580, 20690, 20913, 20529, 20116, 20182, 20276, 20371, 20025, 19942, 20578, 20561, 20181, 19974, 20190, 19301, 19851, 18651, 21292, 10450, 0, 8387, 14795, 14974, 18044, 17129, 17258, 16710, 17052, 17105, 17046, 17164, 16940, 17349, 16537, 19154, 21573, 21070, 21867, 21956, 22189, 22139, 21849, 21794, 21622, 21928, 20682, 19483, 19554, 20470, 21744, 21173, 20648, 20443, 20500, 20504, 20881, 21171, 21439, 21460, 21629, 21758, 21752, 21725, 21773, 21524, 20695, 20197, 20411, 20287, 19978, 19915, 19991, 20078, 20072, 20035, 20126, 19945, 20323, 18962, 16804, 16624, 17099, 17240, 17581, 18625, 19031, 19336, 20799, 21911, 21947, 22053, 22097, 21606, 20997, 21166, 21470, 21539, 21431, 20965, 20865, 21211, 21313, 21589, 21649, 21644, 21545, 21321, 21385, 21487, 21683, 21826, 21963, 22257, 22196, 22095, 22219, 22236, 22321, 22120, 22513, 21781, 23238, 18559, 14612, 16912, 16117, 17048, 16747, 16700, 16624, 16216, 16396, 16627, 16881, 17072, 17732, 18195, 18383, 19353, 20243, 20011, 20075, 20306, 20024, 20054, 19407, 20769, 18263, 21821, 6732, 5637, 20991, 18266, 21162, 20567, 21038, 20991, 20975, 20969, 21011, 20883, 21010, 20813, 21146, 20556, 21745, 17400, 10740, 11680, 6702, 347, 5143, 8732, 8382, 8850, 8285, 8936, 12324, 13548, 16337, 6954, 0, 825, 0, 141, 65, 0, 1236, 1244, 0, 116, 37, 0, 477, 0, 4324, 11488, 12112, 11056, 10902, 14096, 15080, 17043, 18406, 18563, 18548, 18578, 18503, 18661, 18335, 19347, 20183, 20549, 19087, 17107, 17984, 18193, 14932, 4866, 0, 423, 1283, 3416, 4621, 6377, 7433, 7665, 9451, 15571, 6142, 0, 0, 6275, 20245, 11453, 0, 11283, 18700, 22367, 30451, 19147, 17199, 9437, 0, 552, 0, 167, 0, 81, 0, 283, 0, 1004, 0, 8219, 19347, 16859, 18480, 17496, 17807, 17541, 18549, 18670, 17387, 16827, 18401, 18930, 17933, 17893, 18406, 16683, 10993, 9349, 9405, 9037, 9035, 9636, 11960, 5196, 2312, 2269, 0, 697, 0, 3797, 13811, 17782, 18587, 18432, 18468, 18067, 10176, 5634, 6934, 6140, 6862, 5931, 7488, 3478, 5381, 11424, 11819, 10721, 9384, 13107, 13889, 14262, 15543, 15850, 14532, 14301, 14662, 15205, 15710, 16123, 16986, 18263, 19137, 19605, 19278, 19205, 19187, 18839, 18711, 17714, 17969, 15243, 10637, 7854, 13974, 12516, 9856, 15973, 13373, 12489, 11099, 9381, 10064, 9503, 10173, 9139, 11079, 4846, 0, 466, 0, 0, 2513, 9456, 12894, 12167, 10325, 11462, 13897, 15088, 14491, 14448, 13502, 11659, 11590, 12333, 12183, 14035, 14513, 18361, 9540, 9914, 10909, 7145, 16865, 18166, 19025, 18663, 18423, 18502, 18445, 18711, 15358, 14655, 17264, 16948, 17203, 17069, 17121, 17126, 17066, 17266, 17293, 17108, 17186, 17757, 18766, 19108, 19823, 20096, 17651, 18447, 13418, 9230, 11720, 13317, 15532, 15307, 16188, 16000, 14277, 13477, 13529, 13740, 14128, 14051, 15230, 16357, 16100, 15711, 15807, 15524, 14087, 13674, 14164, 13613, 13771, 14454, 14524, 14737, 14607, 14765, 14514, 14957, 14084, 16881, 19335, 18753, 19181, 19244, 18405, 19180, 18293, 19146, 20328, 17541, 17699, 17021, 17534, 17510, 17908, 19256, 20078, 19742, 19162, 17377, 15528, 15228, 15707, 15293, 15131, 15365, 14854, 15746, 16536, 17024, 17809, 18407, 18417, 18102, 17351, 15950, 13696, 13024, 13132, 13139, 13035, 13276, 12764, 14499, 16470, 16636, 17604, 18029, 18827, 19310, 16697, 14922, 14651, 16068, 17356, 16535, 15300, 13791, 14843, 15584, 14211, 14414, 16108, 17938, 17299, 17578, 19336, 19353, 19237, 19714, 17065, 11791, 10553, 11630, 11948, 10971, 12469, 15150, 8344, 3301, 1959, 0, 562, 0, 1027, 0, 7609, 16609, 12403, 13031, 12589, 12640, 12302, 12210, 14614, 16929, 18221, 18172, 12647, 4619, 1288, 1450, 1888, 5318, 7355, 6560, 8164, 9548, 13723, 10778, 0, 2843, 2964, 0, 2701, 5398, 2858, 1881, 1891, 354, 0, 13, 0, 0, 0, 0, 1, 0, 24, 0, 978, 6735, 11321, 5118, 2464, 2644, 5853, 10723, 9729, 11008, 11302, 11305, 11554, 11040, 12110, 12825, 12874, 5651, 390, 845, 0, 0, 875, 2407, 1491, 5147, 8195, 8642, 8817, 9341, 11349, 11243, 12315, 8983, 21695, 32894, 30582, 32634, 31099, 31859, 30794, 32512, 29464, 35497, 15709, 0, 1969, 0, 647, 0, 605, 117, 2173, 4116, 7384, 10366, 10465, 6940, 3035, 4431, 2532, 7987, 12933, 12206, 13694, 13148, 13197, 13175, 13792, 10477, 7108, 9225, 9810, 10317, 10918, 10231, 11126, 10706, 11538, 13604, 14200, 14150, 14068, 14357, 14706, 13755, 15635, 11881, 23428, 26446, 4339, 0, 74, 0, 0, 163, 0, 1402, 2702, 6741, 9234, 4544, 7943, 10911, 10240, 10466, 10733, 10139, 10769, 7127, 3886, 5214, 9358, 10170, 14618, 16266, 12148, 14226, 13401, 14059, 13381, 15603, 18922, 16007, 14413, 15228, 14894, 15071, 14981, 15021, 15008, 14990, 15314, 16499, 13800, 12225, 11622, 10721, 10499, 10643, 4300, 0, 732, 0, 1675, 2616, 6540, 10841, 9383, 10043, 10610, 11064, 11650, 12215, 12118, 11822, 11567, 11219, 11000, 10634, 10737, 10437, 12282, 8017, 3551, 5713, 8064, 11100, 12729, 13554, 13505, 13509, 13575, 13419, 13726, 13084, 15335, 18458, 18190, 17109, 18117, 18975, 18580, 20357, 20146, 20771, 17559, 14962, 16292, 15480, 15777, 15815, 15717, 7905, 3712, 4693, 3841, 3719, 7340, 11570, 11098, 11615, 11285, 11375, 11346, 11194, 11200, 11036, 11282, 10897, 11883, 7786, 3297, 4647, 4746, 4756, 4883, 4547, 5215, 3862, 8216, 12212, 11686, 12847, 17164, 21902, 21624, 22574, 20193, 17530, 20299, 20439, 18943, 19340, 18738, 19145, 18239, 20541, 21322, 21452, 18494, 14520, 15680, 14031, 13621, 14501, 12656, 10854, 11034, 10969, 11104, 11503, 11799, 11719, 11632, 11262, 11130, 11204, 11167, 11179, 11186, 11157, 11219, 11092, 11483, 11730, 11694, 12070, 12136, 12181, 12125, 12503, 12471, 12335, 12599, 12312, 12667, 13164, 14715, 15122, 13829, 13593, 14105, 14942, 18723, 17343, 14784, 15785, 14250, 13575, 11395, 15396, 9079, 7863, 13226, 11250, 14875, 8987, 5374, 6590, 5168, 6423, 7212, 7141, 6903, 7557, 6210, 8878, 1846, 4590, 5632, 0, 9234, 11208, 11821, 11643, 11806, 11896, 11852, 12200, 12121, 12032, 12004, 11898, 12289, 11702, 13033, 10078, 8285, 8754, 7797, 8853, 7417, 8565, 10130, 10694, 11504, 11389, 12865, 12996, 12737, 13949, 14109, 12962, 14177, 8667, 3487, 5099, 4201, 4855, 4197, 5178, 2265, 0, 277, 0, 35, 52, 0, 329, 0, 2179, 2950, 4494, 8767, 2919, 1119, 7348, 10999, 11466, 11714, 11976, 12085, 12192, 11891, 12287, 11547, 9126, 11212, 5407, 0, 4589, 9529, 9951, 10319, 10314, 8198, 9226, 11847, 12931, 14700, 13914, 14626, 13724, 15126, 12476, 21890, 34809, 24729, 25422, 11226, 0, 1425, 0, 399, 0, 16, 71, 0, 662, 467, 605, 3730, 4757, 6368, 10129, 12664, 9470, 6270, 4927, 7415, 9163, 9992, 12990, 12054, 12956, 12111, 14572, 17737, 14342, 10425, 10130, 11770, 11701, 11711, 11596, 11849, 11320, 12351, 10369, 15176, 11704, 18380, 32196, 31045, 32057, 32653, 28658, 24576, 20061, 11319, 3490, 0, 205, 116, 0, 2713, 7120, 8553, 12358, 10148, 9015, 12267, 13438, 13133, 12980, 13196, 12905, 11502, 9388, 7697, 8689, 12202, 17768, 20558, 20746, 19605, 18161, 18568, 18358, 18472, 18399, 18458, 18400, 18173, 15544, 14512, 15124, 14615, 16064, 16738, 17264, 17741, 18032, 15108, 12894, 11880, 10767, 11668, 11655, 11488, 10541, 11943, 4975, 0, 2991, 8670, 12146, 12231, 12771, 13458, 13754, 13953, 13862, 14064, 13776, 13659, 13285, 12345, 11382, 9783, 10905, 12308, 11806, 12191, 11744, 12421, 11156, 15274, 19785, 19238, 19911, 19747, 19650, 20029, 19636, 19214, 20317, 20237, 20239, 20200, 19697, 19805, 20120, 19954, 20098, 19035, 19373, 17116, 14493, 15335, 14852, 15294, 12257, 9499, 8211, 6845, 8302, 11752, 13507, 13377, 13765, 13336, 13172, 13132, 13152, 12974, 13110, 12901, 13263, 12608, 13910, 9604, 5062, 6477, 6502, 8623, 10928, 12363, 11808, 12542, 11667, 15199, 19196, 19087, 20558, 20201, 20533, 20782, 20590, 21105, 21003, 20442, 19799, 19292, 19494, 19321, 20176, 20243, 19127, 18788, 15422, 13530, 13742, 13620, 13730, 13393, 13428, 13124, 13190, 13015, 13165, 12944, 13322, 12650, 13957, 9863, 8216, 15498, 13341, 7695, 7896, 10912, 12143, 11648, 12190, 12805, 12764, 13027, 13077, 12835, 12799, 12564, 12815, 12524, 14273, 17962, 21896, 19711, 16235, 15572, 13121, 13958, 14954, 16906, 18165, 17560, 17377, 17363, 16968, 16710, 17967, 16788, 15628, 15994, 15923, 15759, 16227, 15285, 17183, 11031, 5259, 7484, 5464, 8146, 2219, 2816, 11357, 13246, 15113, 15044, 15141, 13178, 12390, 12850, 12351, 13163, 11017, 8599, 9613, 9304, 11243, 12989, 13311, 13377, 13539, 12332, 10590, 11126, 10767, 10619, 8627, 8976, 10741, 10984, 11680, 11061, 12112, 13109, 12621, 13189, 12319, 13933, 8718, 3387, 5708, 3068, 4126, 2258, 0, 311, 0, 111, 0, 158, 0, 557, 0, 3264, 2305, 6549, 13692, 13061, 13938, 13175, 9718, 8796, 13434, 13307, 14141, 13296, 13785, 12732, 15010, 14362, 10964, 9758, 11599, 4839, 214, 7391, 9707, 10795, 10529, 10473, 10843, 9940, 13032, 16298, 15512, 10955, 17515, 24063, 23535, 28255, 26738, 22240, 22965, 10235, 2311, 7121, 1350, 0, 24, 0, 6, 1, 0, 66, 159, 3959, 7647, 6144, 10033, 10983, 6680, 9314, 11100, 12164, 15100, 17423, 19286, 19268, 19327, 19174, 19436, 20069, 19693, 20156, 19414, 20831, 16163, 10867, 11807, 12419, 13968, 15200, 15159, 17655, 11362, 17135, 30766, 31107, 31728, 32033, 27922, 25560, 22107, 11086, 7147, 8238, 3474, 0, 662, 0, 2880, 8868, 7406, 6644, 6594, 9612, 13326, 12846, 13845, 11839, 8289, 7164, 7623, 6255, 10276, 13757, 12876, 13063, 13409, 12309, 16241, 19609, 18242, 19739, 19116, 18338, 18771, 16588, 15506, 15442, 15451, 15744, 15612, 18408, 17866, 18201, 16337, 13692, 12689, 11333, 11882, 12434, 12208, 12945, 11590, 11538, 5613, 0, 4732, 11148, 11914, 13024, 13723, 13749, 14084, 14188, 14011, 13972, 13989, 13991, 13970, 14023, 13913, 14118, 13789, 15641, 16771, 17209, 18035, 17910, 18394, 18391, 19312, 19960, 20125, 20207, 21009, 20450, 19675, 19932, 20499, 20507, 19447, 19529, 20027, 20455, 20625, 20783, 18747, 18596, 17018, 14567, 15135, 15107, 15157, 14848, 12478, 7798, 7643, 8884, 11427, 13665, 13261, 13503, 13379, 13418, 13462, 13317, 13596, 12897, 13960, 11342, 11299, 16163, 13967, 14706, 10063, 5814, 7899, 10594, 13284, 12773, 12889, 14018, 18194, 19139, 18261, 19639, 20040, 20046, 20542, 20040, 19776, 20094, 20348, 20386, 20005, 19986, 19794, 19855, 19658, 20017, 18482, 19208, 16046, 12518, 13951, 13301, 13603, 13531, 13407, 13776, 12694, 12843, 11865, 11865, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17241, 16334, 16583, 16526, 16422, 16727, 16040, 18319, 20475, 20164, 21073, 21068, 21779, 21513, 22445, 23408, 23735, 24078, 24268, 25499, 23971, 22459, 21214, 19974, 19781, 19685, 19590, 19387, 20302, 22164, 21817, 21821, 22778, 23095, 23983, 23943, 24051, 23974, 24039, 23657, 24953, 25908, 26051, 26141, 26467, 27183, 26912, 27103, 26901, 27193, 26654, 28376, 30028, 29480, 29625, 29789, 29731, 29524, 29865, 30000, 30262, 30393, 30348, 30591, 31118, 31483, 31745, 32505, 31452, 33356, 30769, 36798, 16355, 0, 2360, 0, 1001, 374, 380, 1435, 15, 2643, 0, 16164, 36750, 29654, 31691, 29966, 30130, 29252, 29871, 28985, 30536, 27684, 33365, 14760, 0, 1833, 0, 524, 0, 106, 0, 0, 0, 0, 0, 1, 0, 6, 0, 19, 0, 165, 491, 283, 260, 0, 1000, 1642, 1275, 1030, 0, 54, 0, 14, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 39, 106, 1966, 2576, 1961, 5723, 6834, 12631, 17657, 18508, 19656, 19363, 21374, 21871, 22865, 23180, 23449, 23722, 24103, 24566, 24778, 24922, 24861, 24930, 24817, 25017, 24678, 25091, 20768, 17480, 18695, 15964, 12874, 14683, 8265, 2857, 5004, 4141, 4544, 4130, 4090, 3955, 3833, 3705, 3773, 4061, 4363, 4488, 4646, 4514, 4663, 5056, 5138, 5072, 5032, 4845, 4708, 4420, 4128, 4057, 3274, 897, 0, 83, 0, 53, 0, 149, 0, 500, 0, 4282, 11034, 10782, 13670, 14853, 14905, 17353, 22048, 24521, 24108, 24033, 25366, 25259, 25830, 26262, 24435, 26360, 27438, 27141, 22598, 21455, 19261, 16537, 12529, 1910, 0, 46, 0, 18, 0, 0, 0, 0, 7, 0, 915, 7136, 12250, 12487, 12645, 12480, 12676, 12353, 13424, 14799, 14312, 16949, 19027, 19437, 20637, 21093, 24105, 27050, 28186, 28612, 29039, 28577, 28767, 28128, 29035, 25691, 22680, 20562, 8689, 3297, 3543, 2526, 2467, 2275, 2454, 2791, 2908, 1664, 179, 77, 0, 16, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 30, 0, 120, 0, 840, 1723, 3253, 2095, 0, 1699, 4466, 6376, 7265, 7521, 8641, 8591, 8407, 6145, 5369, 5853, 3224, 765, 0, 68, 0, 15, 0, 2, 0, 0, 0, 1, 0, 5, 0, 20, 0, 162, 150, 0, 22, 0, 6, 0, 5, 0, 19, 0, 77, 0, 823, 2898, 3925, 2875, 5420, 10145, 12156, 14211, 15394, 16839, 18371, 20209, 21141, 21813, 24004, 24401, 23260, 24989, 25994, 25921, 27472, 28401, 29859, 30070, 29564, 29770, 29622, 29775, 29565, 29960, 28660, 27059, 26158, 23773, 20779, 19778, 12268, 1662, 0, 20, 0, 3, 0, 0, 3, 0, 243, 1341, 1716, 1974, 857, 0, 104, 0, 30, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 10, 0, 39, 0, 332, 900, 2110, 7163, 11893, 15458, 17302, 16944, 17072, 17052, 16953, 17205, 16704, 17735, 14065, 8718, 8780, 8132, 6066, 6297, 6425, 6122, 7211, 7224, 6575, 6548, 4983, 1301, 117, 0, 4, 0, 0, 0, 0, 0, 0, 14, 0, 68, 0, 229, 0, 2190, 6851, 7346, 9632, 9984, 10153, 11666, 10777, 10945, 11191, 11184, 11070, 11347, 10794, 11931, 8145, 4111, 5029, 4530, 4615, 4264, 3754, 1406, 0, 42, 0, 10, 0, 0, 2, 0, 0, 514, 5761, 13362, 16248, 17570, 18993, 19403, 19892, 20320, 20946, 21159, 21257, 21469, 21233, 20934, 21049, 20745, 20443, 19456, 18823, 18523, 17903, 18226, 17850, 18451, 17385, 19469, 13052, 7696, 4085, 0, 579, 0, 152, 0, 25, 0, 9, 0, 42, 0, 324, 814, 2025, 3110, 3961, 5332, 6578, 8761, 9028, 9207, 10952, 14444, 19554, 22008, 22815, 22952, 23245, 23846, 24328, 23830, 22741, 23042, 23118, 22723, 22517, 22594, 22514, 22640, 22429, 22840, 21468, 19690, 18815, 14728, 10335, 4849, 479, 0, 0, 0, 19, 0, 62, 304, 4991, 8755, 7876, 10234, 12248, 12618, 12410, 11954, 11142, 12365, 14327, 13789, 12822, 12029, 11328, 10016, 7792, 5182, 4366, 2463, 4066, 6907, 7299, 7711, 7296, 7495, 7351, 7510, 7268, 7720, 6331, 5522, 6498, 6168, 5173, 4346, 5122, 6502, 6729, 7069, 9176, 9912, 10914, 12138, 11165, 8408, 7104, 6657, 1974, 0, 191, 0, 56, 0, 10, 0, 0, 18, 0, 66, 0, 615, 1862, 2208, 1304, 776, 622, 464, 896, 630, 954, 439, 1340, 0, 5416, 11480, 9179, 10404, 10951, 11059, 10174, 11857, 13147, 14616, 16045, 16048, 16350, 16284, 16660, 16727, 16428, 16100, 16336, 16332, 16170, 15522, 15995, 14022, 12908, 7272, 304, 148, 0, 47, 19, 398, 550, 716, 900, 944, 372, 0, 54, 0, 63, 0, 184, 0, 1497, 3692, 3848, 4740, 4690, 4757, 4153, 2570, 588, 0, 49, 0, 13, 0, 0, 0, 0, 0, 128, 1143, 2406, 3465, 5234, 6109, 7476, 9356, 10605, 11169, 11721, 12948, 13490, 14568, 15701, 17994, 20073, 24500, 28042, 28770, 29656, 29342, 29498, 29429, 29448, 29466, 29373, 29201, 28496, 26475, 23011, 16251, 10958, 9673, 9303, 10252, 7227, 4828, 4364, 8129, 8639, 4829, 4744, 3835, 4081, 3610, 3300, 2809, 2770, 2860, 2412, 1970, 1472, 0, 2337, 5832, 7064, 10433, 12085, 13063, 13589, 13872, 13858, 14127, 14416, 14195, 14549, 13915, 15067, 12776, 20365, 28523, 26633, 27922, 27363, 28055, 25918, 23295, 11350, 2882, 4215, 3880, 4529, 4348, 4134, 3105, 2005, 1240, 1145, 1106, 740, 745, 1626, 1655, 1878, 1796, 532, 0, 85, 0, 143, 0, 1427, 5624, 8450, 10280, 11490, 12562, 12907, 12815, 12879, 12803, 12918, 12693, 13391, 14002, 14299, 14314, 16479, 18449, 18834, 19452, 19908, 21944, 20766, 17846, 15763, 8227, 3719, 4472, 4111, 4870, 5731, 6505, 6854, 6718, 7348, 7342, 8008, 9473, 9411, 10046, 10384, 10772, 11424, 11787, 11867, 12002, 12014, 11927, 12013, 12165, 12264, 12160, 12351, 12000, 12644, 11352, 15725, 20898, 19579, 19377, 17892, 16272, 15883, 16610, 16703, 17143, 18892, 20195, 22724, 25255, 26292, 27536, 27885, 28249, 28424, 28322, 28205, 28260, 28535, 28883, 28883, 28974, 29444, 28676, 28071, 23744, 16266, 13636, 13495, 12233, 13183, 7223, 1042, 3557, 4412, 4235, 4450, 4078, 4732, 3460, 7600, 11940, 11074, 12980, 14235, 17498, 21174, 23703, 25081, 25277, 25613, 25866, 25755, 25897, 25762, 24717, 23983, 24181, 23994, 24431, 25561, 25863, 25700, 25698, 26018, 25723, 25908, 25056, 22939, 17727, 10490, 2710, 0, 258, 0, 68, 0, 12, 0, 0, 5, 0, 32, 0, 110, 0, 1652, 5150, 7791, 9872, 10060, 13567, 19945, 24044, 25662, 26517, 27039, 27550, 28162, 28295, 28608, 28917, 28781, 28816, 28528, 28021, 28124, 27999, 28655, 29074, 29466, 30682, 31361, 31374, 31516, 30988, 32568, 28989, 36127, 16372, 0, 2830, 0, 1958, 0, 2842, 0, 15277, 31268, 25776, 19372, 7405, 8597, 7464, 9179, 10745, 11243, 11946, 12325, 12582, 12887, 12969, 13164, 13358, 13406, 13467, 13556, 13514, 13451, 13552, 13361, 13160, 13046, 12971, 13526, 14085, 13715, 13446, 12956, 13726, 13420, 14683, 18518, 19716, 20751, 18794, 17436, 17484, 18038, 16707, 19545, 10158, 1321, 3965, 1380, 2073, 1599, 1280, 1350, 3406, 5947, 3582, 3598, 2741, 315, 1738, 2627, 4584, 6207, 7781, 9321, 10107, 10268, 10502, 10543, 10569, 10572, 13105, 19476, 23548, 24256, 24693, 24528, 24308, 24469, 23176, 21916, 22340, 23008, 23395, 23211, 23435, 23072, 23766, 22329, 26951, 30772, 31937, 29849, 35967, 16052, 0, 2647, 0, 1927, 1331, 1720, 1692, 1418, 2373, 975, 3623, 0, 14820, 31306, 25003, 19923, 13864, 16453, 13495, 13806, 14668, 15170, 15288, 15345, 15447, 15400, 15267, 15296, 15309, 15283, 15321, 15343, 15360, 15341, 15375, 15309, 15436, 15171, 16121, 18472, 22957, 26671, 27151, 27753, 28174, 28430, 28505, 28782, 28790, 29393, 30198, 30802, 31631, 31910, 31461, 31887, 30594, 30567, 15906, 391, 387, 0, 109, 0, 84, 1785, 4654, 5700, 7417, 5634, 2298, 4627, 7455, 8234, 8637, 9196, 9395, 9307, 9425, 9226, 9586, 8864, 11231, 13675, 12988, 12432, 11815, 11782, 11860, 14174, 16427, 18074, 20863, 22752, 23111, 24367, 24926, 25283, 25804, 26619, 28127, 27757, 28242, 28778, 28511, 28761, 28731, 28781, 28892, 26927, 25377, 24479, 22974, 16937, 12897, 13996, 13588, 13919, 13750, 13786, 13775, 13755, 13810, 13711, 13886, 13535, 14799, 16851, 17156, 18724, 19540, 20683, 22568, 23902, 25168, 24776, 24445, 24297, 25994, 27664, 26762, 26721, 27523, 28456, 28866, 28289, 28125, 28621, 27369, 27312, 22612, 17676, 13809, 9448, 10826, 8592, 7280, 7083, 6119, 6197, 5981, 6674, 6822, 7086, 7297, 7194, 7317, 7124, 7460, 6801, 8964, 11241, 10717, 11114, 11162, 11400, 11161, 11470, 11370, 13086, 17292, 19482, 21454, 21274, 20606, 17009, 14069, 15174, 14834, 15104, 15004, 14675, 13988, 13406, 12819, 12531, 11911, 10727, 10009, 9489, 8544, 9073, 10321, 10952, 11801, 12327, 12656, 12591, 12452, 12510, 12457, 12528, 12410, 12638, 11903, 11211, 11391, 11448, 11540, 11408, 10611, 9961, 11130, 10716, 11556, 9749, 8080, 8589, 9334, 10450, 9285, 9629, 9689, 9936, 10281, 11182, 12524, 12524, 12553, 13047, 13114, 13093, 12958, 12884, 12909, 12325, 11869, 11194, 10395, 9904, 10167, 11657, 12150, 12012, 12143, 11953, 12273, 11657, 13646, 15570, 14897, 15258, 15131, 15278, 15032, 14999, 14995, 14658, 14493, 14087, 14078, 13064, 11622, 11789, 11259, 10644, 11105, 11461, 12346, 13073, 12963, 13228, 12534, 13273, 15926, 16205, 16143, 17045, 17609, 18891, 20623, 22219, 23041, 23373, 23903, 22571, 21559, 21995, 21499, 22270, 20928, 23552, 15026, 6544, 8792, 8332, 10167, 10796, 12625, 13536, 14103, 14384, 14567, 14847, 14993, 15158, 14983, 15339, 15170, 16184, 17654, 17478, 18551, 19148, 20117, 21959, 23136, 23161, 23844, 23725, 26050, 28937, 29061, 30131, 30631, 31038, 31311, 31466, 31858, 32240, 32099, 32462, 31767, 32997, 30828, 35243, 18315, 0, 18268, 35279, 29139, 27454, 17016, 12972, 13252, 13004, 12988, 12703, 12528, 12470, 12418, 12352, 12481, 12011, 11272, 11179, 11205, 10653, 10196, 10063, 9554, 8821, 8942, 8571, 7555, 7365, 7396, 4854, 2997, 3447, 3431, 3522, 3338, 3525, 3613, 3633, 3547, 3733, 3380, 4091, 1760, 0, 2319, 2658, 2104, 2629, 1160, 0, 111, 0, 0, 170, 0, 1730, 4608, 2679, 781, 109, 0, 11, 0, 0, 1, 0, 19, 0, 350, 2033, 4072, 5589, 7336, 9744, 11028, 11767, 12187, 12035, 12154, 12346, 12507, 12410, 12545, 12310, 12732, 11891, 14684, 17937, 18275, 19616, 20264, 21460, 22206, 22424, 22404, 21864, 21673, 21966, 21569, 22419, 22047, 22224, 22652, 22728, 22294, 20508, 21520, 16884, 13142, 14583, 14546, 14822, 14851, 15306, 15513, 15721, 15962, 16260, 16367, 16398, 16629, 16726, 16844, 16897, 16845, 16874, 16845, 16886, 16817, 16955, 16490, 15863, 15643, 15421, 14856, 14753, 13508, 11410, 7111, 7162, 11970, 17294, 21443, 22264, 23338, 23937, 23411, 23817, 19669, 15009, 16881, 16192, 10659, 4552, 6069, 3088, 0, 400, 0, 113, 0, 23, 0, 0, 0, 0, 0, 0, 45, 0, 222, 0, 776, 0, 6229, 13862, 10856, 11747, 11165, 11376, 11229, 11855, 11993, 12020, 12586, 12915, 13335, 13358, 14103, 14715, 13990, 15111, 19455, 22420, 23756, 25294, 25119, 26204, 23403, 20018, 15555, 11816, 12800, 12529, 12718, 12359, 11747, 11042, 10391, 9809, 8691, 7859, 7847, 7820, 7835, 7831, 7827, 7841, 7797, 7865, 8380, 8992, 9658, 10104, 9933, 9459, 8325, 7293, 7204, 7252, 7814, 8361, 8832, 9338, 9132, 9167, 8212, 7231, 6327, 1812, 0, 95, 54, 0, 892, 1454, 7257, 12894, 13710, 11078, 7115, 5951, 3570, 4807, 5757, 5805, 6028, 5802, 6148, 5558, 6708, 2966, 0, 386, 0, 193, 0, 328, 0, 2606, 6533, 6040, 7474, 8834, 9994, 11010, 10606, 10004, 9751, 8877, 8170, 7144, 6800, 6750, 6241, 5912, 5615, 5495, 5418, 5511, 1788, 504, 6221, 8377, 13877, 19441, 21469, 24388, 25161, 26177, 26719, 26167, 27120, 25400, 28842, 16881, 189, 537, 0, 172, 0, 20, 0, 0, 0, 0, 0, 0, 9, 0, 23, 228, 3041, 5409, 5683, 6320, 7341, 8363, 8649, 9005, 9374, 9550, 9779, 8319, 6525, 6959, 2507, 0, 278, 0, 81, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 96, 1228, 4527, 6406, 7251, 8871, 9618, 10273, 10405, 10837, 10428, 9502, 8989, 7643, 6916, 6986, 6840, 7079, 6666, 7470, 4788, 1984, 4111, 3690, 3056, 1149, 0, 1534, 3096, 3256, 5550, 10515, 13795, 15575, 13597, 8865, 7666, 8066, 7708, 7893, 8187, 8556, 8479, 8355, 8617, 8791, 8506, 8913, 9488, 9830, 10047, 10473, 11693, 12045, 11987, 12186, 12741, 13440, 13484, 13504, 13483, 13508, 13469, 13548, 13253, 12746, 12678, 12376, 11959, 11726, 10622, 9810, 9264, 7332, 6398, 6417, 6368, 6581, 6850, 6610, 7842, 8612, 9355, 12999, 15912, 18834, 20579, 17432, 8312, 961, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 104, 0, 367, 0, 3027, 7390, 7729, 9805, 9976, 10050, 10290, 10710, 10987, 11343, 11461, 11198, 11094, 10929, 10849, 10118, 9023, 8771, 7332, 5976, 5696, 5882, 5622, 5011, 6288, 7921, 6763, 6856, 8160, 7688, 4943, 2490, 895, 0, 109, 0, 28, 0, 4, 0, 0, 0, 0, 0, 0, 0, 39, 0, 193, 0, 670, 0, 5594, 13649, 12235, 14427, 15057, 16145, 18289, 18532, 20362, 22614, 23932, 25547, 25547, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 4, 0, 30, 0, 1750, 11457, 15601, 10425, 19247, 20278, 14829, 16573, 16287, 17164, 16776, 17572, 17395, 18017, 18822, 19242, 19398, 19321, 19699, 20079, 20227, 20223, 20848, 20140, 21991, 23822, 23320, 24202, 23204, 22879, 22608, 23301, 21938, 24732, 15231, 4220, 7213, 6167, 6403, 6947, 5640, 5181, 2144, 0, 265, 0, 75, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 137, 0, 475, 0, 9116, 9816, 10392, 25377, 27177, 26127, 26529, 26119, 26686, 25781, 27466, 22067, 16764, 18856, 18640, 19445, 19530, 19608, 19828, 20774, 20350, 21599, 24185, 23888, 23699, 22666, 23049, 21889, 26631, 27390, 20593, 21756, 21812, 20103, 18155, 16847, 10066, 4211, 3222, 3319, 1639, 0, 208, 0, 54, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 0, 175, 0, 672, 0, 4831, 7795, 6073, 2098, 8700, 25590, 28032, 29072, 29175, 26524, 22384, 21894, 21731, 20935, 20602, 20386, 19883, 19809, 19524, 19500, 20149, 19721, 23535, 25701, 28668, 33962, 28358, 35869, 16618, 0, 3402, 20, 2246, 326, 2679, 0, 11036, 21062, 13474, 6266, 0, 483, 0, 120, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 149, 0, 575, 0, 4325, 8194, 9310, 5428, 8872, 17988, 24501, 32141, 29554, 29575, 27265, 23892, 22583, 22887, 22739, 22833, 22744, 22866, 22486, 21914, 22088, 21852, 21588, 21608, 21696, 21422, 24155, 24850, 22112, 13037, 4532, 3751, 21064, 29573, 19914, 23458, 26303, 23013, 20597, 7728, 1445, 5166, 4757, 2479, 0, 325, 0, 79, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 150, 0, 594, 0, 3461, 2486, 8708, 23935, 28272, 30969, 30504, 30548, 30103, 30062, 29393, 28370, 30433, 30797, 31678, 29320, 35582, 16929, 0, 1899, 104, 1477, 2350, 3726, 3203, 3932, 2540, 3191, 1523, 3778, 0, 16475, 34822, 28223, 29306, 23976, 24608, 24369, 23963, 25132, 22807, 27479, 12156, 0, 1510, 0, 432, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 563, 4579, 7695, 4018, 8727, 18366, 24099, 30576, 31510, 30873, 29377, 28929, 25134, 21458, 22346, 21571, 21405, 21195, 21154, 21402, 20830, 21944, 19873, 24006, 10556, 0, 2284, 0, 2392, 493, 5184, 0, 17628, 35552, 26204, 27333, 24714, 25121, 18020, 4754, 54, 655, 643, 0, 2493, 7671, 7674, 8230, 8586, 8662, 8967, 8231, 7134, 5923, 5855, 7410, 8110, 8378, 8110, 7458, 7234, 5655, 4606, 4956, 4682, 5010, 4505, 5452, 2406, 0, 299, 0, 85, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 90, 0, 445, 0, 1564, 0, 13114, 32649, 30673, 29158, 25933, 22451, 18352, 19682, 18926, 19737, 20816, 22449, 24945, 29277, 27143, 34838, 15734, 0, 3505, 1298, 4927, 4714, 5135, 4728, 5140, 5780, 5602, 6750, 4311, 7395, 0, 19300, 30215, 18592, 11351, 0, 2936, 434, 1348, 855, 1102, 932, 1151, 510, 0, 63, 0, 18, 0, 15, 0, 59, 0, 200, 0, 1708, 4391, 3603, 3185, 1111, 0, 81, 0, 26, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 112, 0, 404, 0, 3651, 9449, 5639, 0, 7410, 22907, 26119, 24645, 24472, 20779, 18308, 19265, 18840, 19609, 20350, 20679, 21123, 21487, 21346, 21582, 21977, 21936, 21828, 21900, 21711, 21151, 22058, 20241, 23723, 17093, 32599, 13147, 10594, 33716, 20060, 26126, 24231, 24388, 23114, 18402, 15749, 11617, 5805, 5810, 5675, 5786, 5743, 5952, 5570, 6449, 2784, 0, 335, 0, 56, 29, 0, 270, 0, 2157, 4393, 2853, 3163, 1377, 54, 26, 0, 13, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 163, 0, 570, 0, 4577, 10410, 8529, 9657, 8711, 9833, 7967, 13732, 19404, 17886, 18767, 18934, 20007, 20623, 20985, 20997, 21510, 21696, 21319, 21798, 22029, 23805, 25946, 24810, 24740, 23362, 21709, 22112, 19785, 19933, 21028, 22264, 17386, 8263, 6782, 6141, 5663, 5021, 5352, 7640, 8271, 6088, 4774, 4767, 4463, 4500, 4516, 4416, 4638, 4210, 5073, 2244, 0, 278, 0, 79, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 199, 0, 740, 0, 4651, 4412, 5881, 21180, 26125, 21496, 16906, 18239, 17801, 17162, 17448, 18332, 18429, 20686, 21949, 21808, 21799, 21577, 22258, 22362, 21981, 22718, 25183, 27214, 27171, 26014, 25535, 25612, 25645, 25519, 25773, 25292, 26590, 24343, 16168, 19863, 22328, 13504, 7112, 5144, 3047, 292, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 182, 0, 623, 0, 4960, 10302, 5036, 4060, 3487, 1188, 0, 119, 0, 30, 0, 7, 0, 0, 0, 0, 0, 0, 4, 0, 23, 0, 81, 0, 1208, 3312, 4270, 5065, 4266, 2827, 1690, 1233, 1161, 327, 0, 29, 0, 8, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 157, 0, 608, 0, 3729, 3216, 5558, 13727, 17449, 25413, 27887, 29595, 29586, 29484, 28213, 30666, 28152, 34753, 16193, 0, 3095, 0, 1923, 2033, 2201, 2634, 2755, 3128, 3180, 4170, 5246, 5164, 4950, 4771, 2298, 4912, 0, 16971, 35149, 29904, 31988, 31842, 30098, 34878, 17221, 0, 8190, 20148, 9970, 474, 5036, 1076, 0, 41, 0, 27, 0, 18, 0, 32, 0, 116, 0, 763, 763, 0, 116, 0, 32, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 114, 0, 416, 0, 5961, 9871, 11359, 12396, 11756, 7006, 6800, 21583, 26986, 20315, 16957, 18085, 17613, 17664, 18145, 19264, 19087, 19499, 19308, 19451, 19294, 19523, 19086, 20702, 23521, 23165, 25548, 28172, 30767, 29267, 34573, 18260, 0, 19515, 34800, 28460, 27326, 24655, 20214, 13834, 4890, 0, 1087, 367, 726, 504, 367, 116, 213, 277, 108, 0, 12, 0, 7, 0, 22, 0, 77, 0, 627, 1408, 1184, 1270, 1270, 1184, 1408, 627, 0, 77, 0, 22, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 110, 0, 456, 0, 2297, 0, 6341, 17362, 16966, 18210, 18061, 19454, 19465, 20238, 20656, 21782, 22449, 22746, 22984, 22905, 23166, 23378, 23265, 23153, 22503, 22910, 22040, 24662, 26324, 27574, 31528, 32827, 27580, 26096, 15415, 5323, 7816, 5354, 5780, 6024, 6053, 5440, 5535, 5363, 5662, 5128, 6183, 2735, 0, 339, 0, 97, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 59, 0, 245, 0, 2284, 6374, 6088, 166, 9298, 25932, 25855, 25440, 22239, 19376, 20985, 22193, 24578, 26677, 27552, 28260, 28381, 28095, 27701, 28561, 25698, 22953, 23835, 23260, 23826, 23028, 24769, 26606, 34446, 20275, 0, 18203, 31100, 27267, 18563, 5317, 8794, 5220, 3501, 485, 0, 22, 0, 12, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 58, 0, 287, 0, 1006, 0, 8230, 19298, 16822, 18278, 18796, 21132, 21681, 22104, 22000, 22247, 22351, 22254, 21623, 21605, 21295, 20965, 22165, 22398, 24860, 26549, 26438, 35006, 18544, 0, 18600, 33830, 28157, 28691, 25977, 25859, 22691, 12001, 2419, 5790, 3114, 0, 397, 0, 117, 0, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 0, 67, 0, 206, 0, 2221, 6012, 73, 5776, 22957, 26361, 24917, 21511, 19049, 19878, 19624, 20409, 19861, 20250, 21022, 21022, 21113, 21434, 21253, 20946, 21428, 21236, 20780, 21156, 20781, 20830, 21179, 21206, 20921, 21570, 20311, 22862, 14430, 5711, 7985, 6075, 6159, 5787, 5825, 5918, 5078, 3682, 1166, 0, 126, 0, 35, 0, 6, 0, 0, 0, 0, 0, 5, 0, 27, 0, 103, 0, 890, 2483, 2904, 1164, 0, 138, 0, 39, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 117, 0, 492, 0, 3288, 3138, 1184, 0, 11928, 26062, 21239, 23588, 22298, 23039, 22549, 23044, 21788, 20592, 21262, 21525, 21472, 21351, 21648, 21659, 21750, 21632, 21955, 23559, 26375, 25575, 27810, 33274, 29983, 25410, 13313, 3657, 3626, 2507, 2854, 2541, 2166, 1981, 1610, 357, 0, 25, 0, 7, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 100, 0, 361, 0, 3039, 7454, 4898, 1015, 3578, 18973, 21134, 17295, 19293, 18426, 19427, 18947, 18950, 19756, 20738, 20976, 20679, 20514, 20808, 21716, 21680, 21349, 21561, 21639, 21652, 21887, 21786, 27999, 22449, 34718, 11478, 13756, 33133, 16559, 23715, 19695, 22299, 20058, 23119, 14216, 5362, 7080, 6041, 8383, 2780, 0, 295, 0, 94, 0, 21, 0, 0, 5, 0, 24, 0, 86, 0, 606, 838, 0, 46, 0, 13, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 6900, 18120, 21442, 7702, 26514, 20390, 15376, 8258, 3444, 4936, 4162, 4564, 4382, 4410, 4816, 6640, 8402, 10036, 10578, 16472, 29586, 14322, 0, 12190, 24346, 25204, 28404, 28178, 28864, 28220, 30744, 29656, 29554, 27986, 25366, 26530, 30332, 30050, 30130, 31832, 28104, 30612, 32352, 31532, 30054, 31260, 28078, 26370, 31796, 32052, 34508, 35518, 34394, 34904, 34514, 34932, 34344, 35400, 32038, 29070, 31622, 29868, 30798, 30252, 28460, 28968, 27876, 23908, 5272, 13756, 4426, 9860, 5024, 21568, 13610, 13878, 13212, 14630, 18938, 4330, 11506, 3750, 9152, 1796, 8682, 0, 7524, 12488, 14190, 14500, 14216, 6604, 0, 1468, 0, 5522, 11824, 10008, 10848, 10528, 10436, 11088, 8030, 1338, 0, 0, 80, 0, 394, 0, 2694, 2700, 0, 412, 0, 116, 0, 22, 0, 0, 26, 0, 104, 0, 330, 0, 3432, 10604, 5718, 0, 762, 0, 3410, 0, 5776, 724, 11962, 16244, 0, 5016, 5732, 6120, 6114, 5698, 6600, 4896, 9000, 5480, 4358, 9450, 5640, 8076, 12078, 11924, 17400, 21164, 20890, 15782, 15430, 18712, 18516, 24586, 27484, 16208, 14452, 14114, 5788, 1024, 3378, 5000, 0, 3390, 2288, 0, 314, 0, 98, 0, 0, 36, 0, 152, 0, 1240, 2784, 2334, 2518, 2506, 2336, 2810, 1178, 0, 1008, 6988, 4786, 0, 2088, 0, 10152, 11548, 0, 6940, 0, 13696, 14482, 0, 2322, 0, 866, 0, 918, 0, 5262, 5428, 0, 1152, 0, 3284, 7488, 1758, 644, 1192, 0, 214, 0, 60, 0, 0, 90, 0, 464, 0, 1630, 0, 13096, 29334, 24564, 27116, 26092, 24132, 22004, 16944, 11866, 12674, 11534, 12690, 12762, 12004, 14664, 9874, 15138, 21234, 18732, 12848, 11656, 19250, 21796, 28692, 34286, 36464, 36236, 35434, 35906, 34856, 35420, 33240, 31594, 33508, 33346, 31308, 31730, 24150, 17524, 19182, 18910, 18074, 20544, 11450, 744, 5010, 3434, 6012, 316, 14042, 6852, 7096, 10674, 2462, 24676, 8304, 196, 3164, 0, 760, 0, 504, 0, 3670, 10444, 13686, 11918, 5738, 11926, 22924, 25128, 31260, 31440, 24314, 26836, 31502, 22326, 13430, 15202, 15258, 814, 10188, 24982, 20396, 22526, 21722, 21502, 22776, 15558, 7788, 3740, 824, 1556, 358, 9616, 15446, 17248, 17438, 602, 10328, 26260, 27832, 33160, 31000, 31272, 33354, 35968, 33830, 35518, 35372, 33848, 34832, 33038, 33770, 33392, 32172, 29640, 25606, 26514, 28756, 23464, 18704, 18846, 19052, 22498, 24162, 24210, 24222, 24260, 24136, 24396, 24160, 28410, 31464, 30914, 30066, 31378, 31612, 27434, 30848, 29938, 21784, 30562, 19432, 23080, 7644, 11492, 12394, 4046, 8742, 2304, 7122, 94, 7368, 0, 14304, 13018, 0, 3592, 0, 4268, 12082, 15382, 18246, 16354, 4704, 0, 450, 0, 132, 0, 0, 114, 0, 686, 0, 2558, 0, 16606, 14776, 0, 0, 13704, 13444, 0, 0, 16856, 18680, 0, 2892, 0, 908, 0, 660, 0, 2770, 930, 4448, 13616, 9612, 18900, 21264, 16232, 4136, 5822, 27770, 16778, 24978, 23284, 20952, 28126, 3782, 2110, 5718, 4308, 5544, 4040, 6270, 2208, 15188, 23818, 2856, 9854, 30804, 23558, 17770, 26050, 27674, 29942, 28638, 25234, 22180, 19808, 23800, 29668, 29200, 29046, 26608, 22646, 20078, 11030, 2138, 20478, 12568, 0, 0, 6912, 8440, 0, 1316, 0, 340, 0, 64, 0, 0, 0, 0, 0, 38, 0, 134, 0, 394, 0, 4690, 16276, 6758, 0, 2522, 9710, 23082, 6654, 4452, 9168, 0, 5454, 0, 27106, 26718, 0, 4324, 0, 3268, 3628, 0, 9202, 8378, 0, 634, 494, 0, 7626, 7978, 0, 1396, 0, 3836, 4334, 0, 3074, 5874, 4860, 5824, 4470, 6722, 2386, 16304, 29736, 27042, 28634, 25610, 23804, 21886, 27084, 19508, 14314, 16950, 13834, 18830, 17726, 19760, 25264, 21360, 23384, 14876, 18192, 29508, 25186, 26558, 28948, 31590, 33780, 35734, 36444, 35686, 36192, 34764, 32658, 32556, 33480, 32542, 30322, 29158, 21856, 17414, 18772, 17826, 18866, 17332, 20116, 11650, 3528, 2540, 12914, 32022, 14026, 11562, 26384, 10040, 8918, 16950, 6130, 7974, 4678, 7446, 6228, 0, 0, 4388, 16770, 17836, 22120, 14396, 13890, 21772, 23812, 26276, 23294, 29902, 34822, 39262, 27726, 19292, 21602, 20246, 23028, 27856, 23824, 17152, 19260, 18266, 18668, 18718, 18222, 18810, 10634, 7520, 7660, 12032, 20612, 18162, 20746, 19670, 19960, 3412, 9696, 28504, 25218, 30778, 30610, 29628, 32768, 36120, 34906, 35084, 33656, 33568, 35728, 35218, 31050, 31286, 32610, 30824, 25408, 25384, 26170, 24274, 24236, 18422, 22560, 26144, 27204, 28878, 28336, 28494, 28650, 28130, 29236, 26400, 29542, 35052, 33228, 35332, 34946, 33188, 33590, 31272, 31654, 30028, 19158, 10690, 10342, 976, 17968, 15498, 18556, 19910, 0, 17462, 14428, 0, 3668, 5750, 26014, 13882, 0, 2484, 1822, 8508, 15450, 20410, 18200, 4900, 0, 0, 3446, 8502, 6922, 7632, 7346, 7392, 7608, 5154, 0, 9196, 5548, 3160, 3400, 5402, 10882, 0, 25782, 17572, 0, 2430, 0, 616, 0, 0, 1368, 1440, 0, 246, 0, 46, 556, 8078, 21080, 13740, 12396, 21796, 22234, 21974, 30846, 15328, 24232, 19074, 22610, 15730, 6480, 30858, 21882, 25996, 24724, 23724, 27628, 13238, 0, 422, 770, 0, 10478, 17840, 9296, 19904, 28004, 31224, 29704, 29674, 26898, 27610, 29602, 31500, 27464, 25674, 12692, 13392, 19058, 0, 9560, 7684, 0, 3548, 0, 722, 0, 218, 0, 308, 0, 1620, 0, 8802, 8718, 0, 1194, 0, 0, 928, 0, 6898, 7264, 9528, 12014, 64, 150, 516, 0, 5614, 5766, 0, 1368, 0, 2392, 0, 10824, 0, 23786, 26484, 0, 3200, 1094, 4634, 0, 1014, 0, 2014, 1918, 0, 566, 0, 2236, 5048, 5420, 3970, 0, 7706, 13958, 9906, 11350, 11014, 10414, 12160, 8324, 21400, 34382, 24308, 26630, 20136, 12172, 15162, 13324, 17758, 18086, 14814, 11180, 6548, 7170, 4924, 11534, 25342, 9998, 12962, 12130, 8420, 26538, 26120, 31206, 31558, 33364, 36940, 39908, 39066, 39044, 37834, 31760, 30680, 32544, 32124, 30714, 27064, 12444, 5620, 7368, 6486, 7044, 6586, 7124, 5808, 4840, 5398, 5034, 5780, 11352, 32340, 33104, 22958, 26348, 27468, 28400, 26228, 25152, 9212, 4678, 3600, 1024, 1764, 5868, 16298, 18306, 17934, 16626, 1932, 10246, 28472, 29046, 32252, 19490, 17946, 32136, 16534, 11740, 17634, 2898, 4842, 3048, 28, 874, 678, 300, 1420, 0, 6276, 6730, 0, 4378, 2412, 1864, 15054, 20598, 20538, 17244, 11984, 0, 12908, 30096, 29130, 31320, 29470, 34928, 37834, 37262, 39832, 40876, 38068, 35902, 34964, 35228, 36358, 35496, 33068, 29540, 28544, 29156, 28802, 28626, 25598, 26756, 29094, 29666, 30360, 30128, 30198, 30260, 30044, 30482, 29758, 33744, 35118, 32044, 33208, 37012, 32042, 34686, 30180, 32122, 25822, 27858, 10912, 9062, 19214, 0, 1902, 0, 4968, 25616, 18026, 0, 19734, 15690, 0, 3066, 262, 1048, 4504, 15962, 20284, 27186, 38446, 18694, 0, 1480, 0, 440, 0, 86, 0, 0, 0, 0, 0, 2, 0, 0, 164, 0, 896, 0, 3840, 0, 23152, 23050, 0, 3310, 0, 150, 1052, 0, 9984, 10568, 0, 2782, 0, 10804, 25114, 26044, 22142, 18990, 15068, 24438, 29208, 17118, 13310, 18960, 24378, 5390, 3164, 24936, 34176, 31048, 34288, 29338, 38410, 12852, 5934, 9444, 3756, 24988, 22562, 20676, 3614, 17004, 28632, 18872, 28538, 30612, 29672, 29804, 22002, 21148, 14068, 20856, 12230, 20640, 14566, 19098, 21030, 0, 4604, 0, 8848, 722, 13530, 15952, 0, 2530, 0, 604, 0, 432, 0, 64, 0, 156, 0, 596, 0, 3078, 382, 5260, 6870, 0, 2510, 0, 9994, 9582, 0, 1514, 0, 666, 0, 966, 0, 5812, 5812, 0, 886, 0, 248, 0, 48, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 58, 0, 1008, 6280, 14092, 16672, 16412, 15998, 17134, 14660, 23166, 32728, 28544, 32440, 21284, 14112, 13028, 21642, 24806, 9036, 8014, 6610, 6484, 4616, 9806, 13230, 19172, 12256, 2824, 4460, 12294, 24572, 27088, 32714, 32480, 35140, 36596, 38466, 39734, 37466, 32358, 33462, 31418, 32886, 20808, 5034, 7514, 5892, 7036, 6572, 6624, 6932, 6166, 7770, 3460, 5216, 5354, 3488, 2102, 17800, 11384, 0, 0, 13594, 13134, 0, 6886, 0, 8226, 3860, 0, 1454, 10978, 20414, 21564, 17872, 15710, 1746, 9320, 19754, 19846, 22934, 16638, 22504, 28748, 28252, 14752, 11158, 4860, 326, 1444, 0, 1532, 644, 1538, 236, 2504, 0, 11466, 19208, 16424, 12652, 11156, 21202, 18918, 21260, 18942, 7820, 0, 12198, 29430, 29020, 30346, 29958, 33092, 36248, 37206, 38026, 39262, 35544, 34842, 37106, 33750, 34134, 33496, 31650, 30178, 29458, 27750, 25976, 26414, 25830, 26402, 27008, 26830, 26110, 26682, 26374, 26664, 26276, 26916, 25712, 29494, 32228, 29444, 31662, 30614, 23266, 16520, 3388, 25246, 13394, 16178, 10062, 13104, 19102, 0, 7500, 0, 18998, 5362, 8620, 29698, 26792, 28898, 23652, 12574, 10690, 2962, 3982, 14914, 24680, 33830, 31838, 34946, 25884, 9000, 0, 7292, 15044, 11670, 13370, 12086, 13498, 11360, 15356, 4326, 4476, 4546, 790, 0, 18540, 20792, 0, 11254, 23208, 29184, 30408, 12552, 428, 0, 6588, 11128, 0, 21706, 19672, 4082, 21134, 19594, 21810, 22700, 21040, 3692, 7306, 26462, 22052, 19844, 16096, 15866, 28246, 10526, 0, 3954, 0, 822, 0, 346, 0, 564, 0, 5648, 22066, 34450, 33210, 25404, 30690, 30640, 26968, 30104, 24880, 27708, 25078, 26460, 29180, 20158, 21426, 19970, 24908, 7232, 7704, 31184, 13944, 0, 442, 0, 176, 0, 0, 106, 0, 362, 0, 2700, 4586, 0, 7518, 3038, 8006, 22434, 17790, 19676, 19548, 18014, 21978, 8830, 2634, 23802, 7296, 1122, 0, 17708, 11144, 12212, 23638, 0, 20190, 15740, 0, 4392, 0, 15232, 13990, 0, 1612, 614, 1948, 0, 0, 2616, 0, 20202, 18714, 0, 8508, 4398, 0, 374, 0, 0, 1570, 1978, 9512, 16688, 14348, 15784, 14556, 16004, 13592, 21674, 30724, 16462, 16426, 20580, 24130, 27764, 29070, 22960, 12524, 17112, 24146, 16614, 10696, 11728, 20616, 16978, 12822, 20086, 21594, 25386, 20830, 24172, 26624, 25774, 30552, 34334, 35646, 37458, 36896, 34058, 32592, 34958, 32498, 32094, 31768, 28902, 14840, 5824, 8364, 7186, 7644, 7784, 7010, 8074, 1768, 17002, 19118, 0, 984, 0, 3760, 19462, 21896, 4956, 0, 750, 2870, 2322, 0, 1262, 0, 9474, 28838, 26310, 24214, 11440, 0, 10810, 21804, 16578, 21958, 15860, 15462, 23544, 22612, 12552, 17380, 13604, 3308, 25690, 12424, 0, 1228, 0, 0, 1986, 0, 15348, 21706, 13982, 21438, 18988, 25970, 23216, 24602, 19000, 6318, 0, 12140, 25620, 24040, 26942, 28158, 31598, 32102, 31706, 34506, 33932, 31038, 33594, 32530, 29508, 24848, 26982, 27682, 24510, 27210, 25704, 27474, 25360, 23358, 25186, 24858, 23248, 21994, 22776, 22424, 22658, 22438, 22754, 22156, 23948, 24228, 24042, 22340, 25640, 10990, 17178, 10538, 15950, 17220, 0, 2736, 0, 792, 0, 460, 0, 1186, 0, 7776, 7776, 0, 1168, 0, 252, 10, 0, 592, 0, 10050, 22806, 26024, 9296, 0, 0, 6370, 3304, 8594, 24516, 19324, 21516, 21154, 19870, 23572, 10458, 0, 1134, 0, 0, 1196, 6, 4884, 17948, 7108, 0, 738, 0, 0, 380, 1212, 20386, 16978, 18496, 26588, 18570, 29586, 27352, 21926, 25252, 17858, 17614, 14048, 16580, 16604, 24436, 6900, 13964, 14316, 4856, 7158, 8518, 14410, 0, 2040, 0, 0, 1884, 0, 18782, 46138, 23908, 13654, 25908, 32708, 26736, 26796, 27372, 27892, 21886, 21602, 21646, 17242, 19484, 19632, 18820, 25006, 522, 17770, 10840, 14976, 23076, 0, 3858, 0, 1008, 0, 156, 0, 0, 96, 0, 612, 382, 114, 0, 2166, 5118, 4052, 4858, 3910, 5408, 2502, 11380, 14452, 5660, 0, 14516, 8734, 9436, 19552, 0, 21812, 18348, 0, 4716, 0, 12878, 5544, 10512, 14954, 0, 2634, 0, 1170, 0, 5168, 14074, 6154, 0, 5846, 3540, 1536, 1970, 2844, 9288, 7638, 4336, 14084, 13706, 40, 342, 138, 0, 1698, 0, 14204, 31542, 26520, 21478, 19782, 21440, 11070, 6364, 5910, 4254, 10518, 9386, 3152, 5518, 4508, 4880, 4392, 3446, 3512, 12208, 17108, 18728, 24294, 25586, 28920, 32036, 32836, 32796, 29634, 25576, 26798, 28520, 21260, 19584, 18062, 13742, 9468, 5260, 8172, 9716, 9192, 9728, 8942, 10346, 5928, 914, 3494, 2412, 4636, 0, 16508, 11394, 7270, 14104, 7782, 18722, 10308, 18678, 11334, 842, 2504, 16256, 26494, 26096, 22236, 7872, 0, 9300, 17268, 12748, 24534, 18060, 11678, 22426, 9246, 0, 5662, 4038, 0, 1392, 0, 7538, 16806, 14012, 15638, 14426, 15618, 13840, 20278, 30596, 17598, 17476, 26456, 24536, 26172, 14346, 3628, 0, 9760, 23086, 21948, 24914, 24968, 28728, 28654, 29862, 29004, 27764, 27350, 19894, 8972, 7290, 4886, 16740, 25596, 21440, 25394, 23226, 19750, 21906, 14534, 12400, 21328, 16194, 4626, 0, 536, 0, 532, 0, 1424, 0, 11426, 26502, 19918, 23710, 15696, 12164, 24864, 4640, 8084, 3298, 13284, 15096, 0, 0, 15484, 13990, 3750, 13288, 0, 15394, 43244, 18100, 0, 2004, 0, 578, 0, 0, 2434, 17702, 20970, 9682, 1106, 2332, 2954, 0, 464, 0, 120, 0, 10, 30, 0, 200, 0, 832, 0, 5100, 3978, 0, 0, 14054, 48848, 20202, 0, 4240, 0, 16564, 29574, 9860, 4486, 8352, 15490, 28386, 33438, 29404, 31228, 29038, 23982, 22998, 15744, 25778, 7978, 16162, 16288, 16162, 23366, 0, 1534, 214, 0, 11580, 26606, 22514, 23502, 24958, 20466, 30070, 4856, 19838, 26704, 5366, 29986, 26870, 29224, 26928, 22960, 21858, 15856, 7824, 5872, 7090, 5952, 18208, 11130, 12214, 19410, 0, 15720, 13856, 0, 2264, 0, 1904, 798, 42, 0, 1698, 42, 1822, 0, 14364, 14516, 0, 2216, 0, 662, 0, 346, 0, 806, 0, 5180, 4694, 0, 2176, 0, 3574, 16192, 8572, 0, 2068, 0, 3924, 0, 0);

    
    
    -- contador
--    signal r_reg : std_logic_vector(9 downto 0) := "0000000000";
--    signal r_reg : std_logic_vector(10 downto 0) := "00000000000";
    signal r_reg : std_logic_vector(15 downto 0) := "0000000000000000";

begin
-----------------------------------------------------
-- Asignaciones de la arquitectura       
-----------------------------------------------------  
--DEDO_DATA_WR <= x"0000" & tactel(15 downto 0);

--DEDO_ADDR_WR <= "0000" & int_dedo_addr_wr;

DEDO_DATA_WR <= data_tactel_register;
DEDO_ADDR_WR <= address_tactel_register;

-- Salida depuracion r_reg
r_reg_out <= r_reg;

--DEDO_ADDR_WR <= "010" & "0101"; -- SIEMPRE TACTEL 28!!!


ROW_COLUMN <= aux_addr_tactel_register;


-----------------------------------------------------
-- Asignaciones para el bus SPI      
-----------------------------------------------------
ODDR_inst : ODDR
generic map(
        DDR_CLK_EDGE => "OPPOSITE_EDGE",                                    -- "OPPOSITE_EDGE" or "SAME_EDGE"
        INIT => '0',                                                        -- Initial value for Q port ('1' or '0')
        SRTYPE => "SYNC")                                                   -- Reset Type ("ASYNC" or "SYNC")
port map (
        Q => dedo_sclk,                                                     -- 1-bit DDR output
        C => clk,                                                           -- 1-bit clock input
        CE => '1',                                                          -- 1-bit clock enable input
        D1 => '1',                                                          -- 1-bit data input (positive edge)
        D2 => '0',                                                          -- 1-bit data input (negative edge)
        R => '0',                                                           -- 1-bit reset input
        S => '0'                                                            -- 1-bit set input
);

dedo_ss <= int_dedo_ss;
dedo_mosi <= int_dedo_mosi;

-----------------------------------------------------
-- Proceso para dedo_miso que se guarda en tactel                          
-----------------------------------------------------  
process(clk)
begin
    if (clk'event and clk = '1') then
        if state = st5_store_tactels then
            for i in 0 to 30 loop
                tactel(i+1) <= tactel(i);
            end loop;
            tactel(0) <= dedo_miso;
        end if;
    end if;
end process;

-----------------------------------------------------
-- Registro de Operaci�n para el sensor falange0	
-- Carga Paralela Salida Serie							
-----------------------------------------------------	
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st1_idle  then
            reg_command <= "0000000" & dedo_enable; 
        elsif state = st2_send_command then
            reg_command(7 downto 1) <= reg_command(6 downto 0);
        end if;
    end if;
end process;


----------------------------------------------------
-- Registro de estado de la m�quina de estados principal       
-----------------------------------------------------    
SYNC_PROC: process (clk)
begin
    if (clk'event and clk = '1') then
            state <= next_state;
    end if;
end process;


-----------------------------------------------------
-- Salidas de la m�quina de estados principal                     
-----------------------------------------------------    
OUTPUT_DECODE: process (state, reg_command(7), reg_tactel_inicial(7), reg_tactel_final(7))
begin
  case (state) is
        when st1_idle =>
            int_dedo_ss <= '1';
            int_dedo_mosi <= '0';
        when st2_send_command_pause =>
            int_dedo_ss <= '0';
            int_dedo_mosi <= '0';
        when st2_send_command =>
            int_dedo_ss <= '0';
            int_dedo_mosi <= reg_command(7);
        when st3_send_tactel_inicial =>
            int_dedo_ss <= '0';
            int_dedo_mosi <= reg_tactel_inicial(7);
        when st4_send_tactel_final =>
            int_dedo_ss <= '0';
            int_dedo_mosi <= reg_tactel_final(7);
        when st5_store_tactels =>
            int_dedo_ss <= '0';
            int_dedo_mosi <= '0';
        when st7_interno_current_frame_update =>
            int_dedo_ss <= '1';
            int_dedo_mosi <= '0';
        when others =>
            int_dedo_ss <= '1';
            int_dedo_mosi <= '0';
  end case;
end process;


-----------------------------------------------------
-- Pr�ximos estados de la m�quina de estados principal          
-----------------------------------------------------    
NEXT_STATE_DECODE: process (state, byte_counter, row, column, tactel_counter, contador_pausa)
begin
  next_state <= state;
  case (state) is
        when st1_idle =>
             if contador_pausa = "0000101101001101110" then     -- 23150
--             if contador_pausa = "0000110111001011101" then -- 28253 , only for debugging
--            if contador_pausa = "0000000000000100000" then     -- 16 solo para simulacion
                next_state <= st2_send_command_pause;
            end if;
        when st2_send_command_pause =>
            next_state <= st2_send_command;
        when st2_send_command =>
            if byte_counter = "111" then
                next_state <= st3_send_tactel_inicial;
            end if;
        when st3_send_tactel_inicial =>
            if byte_counter = "111" then
                next_state <= st4_send_tactel_final;
            end if;
        when st4_send_tactel_final =>
            if byte_counter = "111" then                    
                next_state <= st5_store_tactels;
            end if;
        when st5_store_tactels =>
--            if row = "111" and column = "1111" and tactel_counter = "11111" then           -- Para leer las dos filas de calibraci�n    
            if row = "100" and column = "1010" and tactel_counter = "11111" then           -- Para leer las dos filas de calibraci�n                  
                next_state <= st7_interno_current_frame_update;
            end if;
        when st7_interno_current_frame_update =>
            next_state <= st1_idle;
        when others =>
        next_state <= st1_idle;
  end case;      
end process;

-----------------------------------------------------
-- Frame Actual (Donde se va a escribir o se est�    
-- escribiendo)                                                
-----------------------------------------------------
process (clk)
begin
    if clk'event and clk='1' then
        if state = st7_interno_current_frame_update and ram_reading = '0' then        -- Cuando se termina la escritura se comprueba si no se est� leyendo
            interno_current_frame <= not interno_current_frame;                               -- y se cambia de bloque      
            contador_one_tactel <= contador_one_tactel + 1;        
            pulso <= '1';
        else 
            pulso <= '0';
        end if;                                                               -- Ojo debe ser s�lo un ciclo
    end if;
end process;

interno_last_frame <= not(interno_current_frame);                             -- Ultimo bloque escrito completo

-----------------------------------------------------
-- Contador de n�mero de ciclos pausa                                     
-----------------------------------------------------    
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st7_interno_current_frame_update then
            contador_pausa <= (others => '0');
        elsif state = st1_idle then
            contador_pausa <= contador_pausa + 1;
        end if;
    end if;
end process;

-----------------------------------------------------
-- Contador para el env�o y recepci�n de bytes        
-----------------------------------------------------
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st2_send_command_pause then
            byte_counter <= "000";
        else
            byte_counter <= byte_counter + 1;
        end if;
    end if;
end process;

-----------------------------------------------------
-- Contador de filas                                            
-----------------------------------------------------    
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st1_idle then
            row <= "000";
--        elsif state = st5_store_tactels and tactel_counter = "11111" and column = "1111" then
        elsif state = st5_store_tactels and tactel_counter = "11111" and column = "1010" then
            row <= row + 1;
        end if;
    end if;
end process;

-----------------------------------------------------
-- Contador de columnas                                        
-----------------------------------------------------    
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st1_idle then
            column <= "0000";
        elsif state = st5_store_tactels and tactel_counter = "11111" then
            column <= column + 1;
        end if;
    end if;
end process;


-----------------------------------------------------
-- Contador para la recepci�n de tactel (4 bytes)    
-----------------------------------------------------    
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st1_idle then
            tactel_counter <= "00000";
        elsif state = st5_store_tactels then
            tactel_counter <= tactel_counter + 1;
        end if;
    end if;
end process;

-----------------------------------------------------
-- Registro para ack_ram_reading                            
-----------------------------------------------------    
process(clk_100)
begin
   if clk_100'event and clk_100='1' then
       if ram_reading = '1' then
           ack_ram_reading <= '1';
       else
           ack_ram_reading <= '0';
       end if;
   end if;
end process;


-----------------------------------------------------
-- int_dedo_addr_wr process                                    
-----------------------------------------------------	
process (clk)
begin
    if (clk'event and clk = '1') then
        int_dedo_addr_wr <= interno_current_frame & row & column;
--        int_dedo_addr_wr <= row & column;
    end if;
end process;	

-----------------------------------------------------
-- Write Enable de la RAM		
-- Escribimos solamente cuando recibimos un 
-- determinado tactel de la matriz, no todos, 
-- ya que el algoritmo por ahora se aplica
-- solamente sobre la secuencia temporal
-- de un solo tactel.
-- En principio voy a poner el tactel (1,5),
-- pero se puede cambiar.							
-----------------------------------------------------
process(clk)
begin
    if (clk'event and clk = '1') then
        if(state = st5_store_tactels and tactel_counter = "11111" and row < "101" and column < "1011") then
            CE_DAT_REG <= '1';                                                  -- Se escribe cuando se han recidido los 32 bits de cada tactel           
        else
            CE_DAT_REG <= '0';
        end if;
    end if;
end process;

-----------------------------------------------------
-- Pasamos la se�al por dos registros - CIRCUITO
-- PULSO						
-----------------------------------------------------
process(clk_100)
begin
    if(clk_100'event and clk_100 = '1') then
        CE_RET_1 <= CE_DAT_REG;    
    end if;
end process;

process(clk_100)
begin
    if(clk_100'event and clk_100 = '1') then
        CE_RET_2 <= CE_RET_1;    
    end if;
end process;

CE_PULSO_100 <= not(CE_RET_1) and CE_RET_2;

-- Maquina de estados FIR - Salida tipo Moore
-- A. Registro de estado de la m�quina de estados FIR
SYNC_PROC_FIR: process (clk_100)
begin
    if (clk_100'event and clk_100 = '1') then
            state_FIR <= next_state_FIR;
    end if;
end process;

-- B. Pr�ximos estados de la m�quina de estados FIR        
NEXT_STATE_DECODE_FIR: process (state_FIR, CE_PULSO_100, t_ready_FIR)
begin
  next_state_FIR <= state_FIR;
  case (state_FIR) is
        when st1_FIR =>
            if CE_PULSO_100 = '1' then   
                next_state_FIR <= st2_FIR;
            end if;
        when st2_FIR =>
            if t_ready_FIR = '1' then   
                next_state_FIR <= st1_FIR;
            end if;
        when others =>
            next_state_FIR <= st1_FIR;
  end case;      
end process;

-- C. Salidas de la m�quina de estados FIR          
OUTPUT_DECODE_FIR: process (state_FIR)
begin
  case (state_FIR) is
        when st1_FIR =>
            t_valid_FIR <= '0';
        when st2_FIR =>
            t_valid_FIR <= '1';
        when others =>
            t_valid_FIR <= '0';
  end case;
end process;



-----------------------------------------------------
-- Registros para el dato y col,fil					
-----------------------------------------------------
--REGISTER_DATA_TACTEL: process(clk_100)
--begin
--    if(clk_100'event and clk_100 = '1') then
--        if(CE_PULSO_100 = '1') then
--            --data_tactel_register <= tactel;
--            data_tactel_register <= std_logic_vector(to_unsigned( reg_datos_debug(to_integer(unsigned(r_reg))) ,32));
--            r_reg <= r_reg + 1;
--        end if;
--    end if;
--end process;

-- THE NEXT PROCESS IS ONLY FOR DEBUGGING
REGISTER_DATA_TACTEL: process(clk_100)
begin
    if(clk_100'event and clk_100 = '1') then
        if(CE_PULSO_100 = '1') then
            data_tactel_register <= std_logic_vector(to_unsigned( reg_datos_debug(to_integer(unsigned(r_reg))) ,32));
        end if;
    end if;
end process;
process(clk)
begin
    if(clk'event and clk = '1') then
        if(state = st7_interno_current_frame_update) then
--            if(r_reg = 32783) then
            if(r_reg = 30734) then    
--            if(r_reg = 16383) then   
                r_reg <= (others => '0');
            else
                r_reg <= r_reg + 1;
            end if;            
        end if;
    end if;
end process;
--process(clk)
--begin
--    if(clk'event and clk = '1') then
--        if(state = st7_interno_current_frame_update) then                
--            r_reg <= r_reg + 1;
--        end if;
--    end if;
--end process;

REGISTER_COL_FIL: process(clk_100)
begin
    if(clk_100'event and clk_100 = '1') then
        if(CE_PULSO_100 = '1') then
            address_tactel_register <= row & column_ret_2;
        end if; 
    end if;
end process;

COLUMN_RET_1_PROCESS: process(clk)
begin
    if(clk'event and clk = '1') then
        column_ret_1 <= column;
    end if;
end process;

COLUMN_RET_2_PROCESS: process(clk)
begin
    if(clk'event and clk = '1') then
        column_ret_2 <= column_ret_1;
    end if;
end process;

REGISTER_ROW_COLUMN_SLOW: process(clk)
begin
    if(clk'event and clk = '1') then
        aux_addr_tactel_register_slow <= row & column;
    end if;
end process;

REGISTER_ROW_COLUMN: process(clk_100)
begin
    if(clk_100'event and clk_100 = '1') then
        aux_addr_tactel_register <= row & column;
    end if;
end process;



-----------------------------------------------------
-- Enable frame number								
-----------------------------------------------------
enable_frame_number <= '1' when state = st7_interno_current_frame_update else '0';


--process(clk)
--begin
--   if (clk'event and clk = '1') then
--       if state = st5_store_tactels then	
--           t_valid_FIR <= '1';
--       end if;
--   end if;
--end process;

-----------------------------------------------------	
-- PROCESO PARA EL START_OUT
-----------------------------------------------------	
div_freq_start: process(clk) 
begin
    if rising_edge(clk) then
        if(contador_start = 4168000) then
            temporal_start <= NOT(temporal_start);
            contador_start <= 0;
        else
            contador_start <= contador_start + 1;
        end if;
    end if;
end process;

START_OUT <= '1' when contador_start < to_integer(unsigned(duty)) else '0';

-----------------------------------------------------	
-- PROCESO PARA EL FRAME_NUMBER STAGE 1
-- STAGE 1: EL FRAME_NUMBER QUE SE PRODUCE AQU�
-- STAGE 2: EL FRAME NUMBER QUE SE PRODUCE EN EL DEDO
-----------------------------------------------------	
frame_number_stage_1: process (clk)
begin
    if (clk'event and clk = '1') then
--        if state = st7_interno_current_frame_update then
        if state = st2_send_command_pause then
            frame_number_stage1 <= frame_number_stage1 + 1;
        end if;
    end if;
end process;
--frame_number <= frame_number_stage1;  

-----------------------------------------------------
-- Registro Frame                                            
-- Carga Serie Salida Paralela                            
-----------------------------------------------------    
process (clk)
begin
    if (clk'event and clk = '1') then
        if state = st2_send_command then
            for i in 0 to 6 loop
                int_frame_number(i+1) <= int_frame_number(i);
            end loop;
            int_frame_number(0) <= dedo_miso;        
        end if;
    end if;
end process;
-- STAGE 2
frame_number <= int_frame_number;  


end Behavioral;